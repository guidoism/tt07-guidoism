/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_guidoism (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // All output pins must be assigned. If not used, assign to 0.
  //assign uo_out  = ui_in + uio_in;  // Example: ou_out is the sum of ui_in and uio_in
  //assign uio_out = 0;
  //assign uio_oe  = 0;

// Generated automatically via PyRTL
// As one initial test of synthesis, map to FPGA with:
//   yosys -p "synth_xilinx -top toplevel" thisfile.v
//
// module toplevel(clk, rst, a, direction, invert, n, shift_in, overflow, s);
//    input clk;
//    input rst;
//   
//    input[63:0] a;
//    input direction;
//    input invert;
//    input[5:0] n;
//    input shift_in;
//    output overflow;
//    output[63:0] s;

   reg [63:0]        a;
   assign a[7:0] = ui_in;
   assign a[63:8] = 0; // We don't have enough pins to set these so they get a zero
   
   wire [5:0]        n;
   wire              direction;
   wire              invert;
   wire              shift_in;
   assign uio_out = 0;
   assign uio_oe = 0;
   assign n[4:0] = uio_in[4:0];
   assign n[5] = 0;
   assign direction = uio_in[5];
   assign invert = uio_in[6];
   assign shift_in = uio_in[7];
   
   wire overflow;
   reg [63:0] s;
   assign uo_out = s[7:0];

    reg[255:0] control_microcode;

    wire const_0_0;
    wire const_1_0;
    wire const_2_0;
    wire const_3_0;
    wire const_4_0;
    wire const_5_0;
    wire const_6_0;
    wire const_7_0;
    wire const_8_0;
    wire const_9_0;
    wire const_10_0;
    wire const_11_0;
    wire const_12_0;
    wire const_13_0;
    wire const_14_0;
    wire const_15_0;
    wire const_16_0;
    wire const_17_0;
    wire const_18_0;
    wire const_19_0;
    wire const_20_0;
    wire const_21_0;
    wire const_22_0;
    wire const_23_0;
    wire const_24_0;
    wire[63:0] reverse_in;
    wire[63:0] reverse_out;
    wire[63:0] shift_1;
    wire[63:0] shift_2;
    wire[63:0] shift_4;
    wire[63:0] shift_8;
    wire[63:0] shift_16;
    wire[63:0] shift_32;
    wire shift_in;
    wire shift_off_1;
    wire[1:0] shift_off_2;
    wire[3:0] shift_off_4;
    wire[7:0] shift_off_8;
    wire[15:0] shift_off_16;
    wire[31:0] shift_off_32;
    wire tmp0;
    wire tmp1;
    wire tmp2;
    wire tmp3;
    wire tmp4;
    wire tmp5;
    wire tmp6;
    wire tmp7;
    wire tmp8;
    wire tmp9;
    wire tmp10;
    wire tmp11;
    wire tmp12;
    wire tmp13;
    wire tmp14;
    wire tmp15;
    wire tmp16;
    wire tmp17;
    wire tmp18;
    wire tmp19;
    wire tmp20;
    wire tmp21;
    wire tmp22;
    wire tmp23;
    wire tmp24;
    wire tmp25;
    wire tmp26;
    wire tmp27;
    wire tmp28;
    wire tmp29;
    wire tmp30;
    wire tmp31;
    wire tmp32;
    wire tmp33;
    wire tmp34;
    wire tmp35;
    wire tmp36;
    wire tmp37;
    wire tmp38;
    wire tmp39;
    wire tmp40;
    wire tmp41;
    wire tmp42;
    wire tmp43;
    wire tmp44;
    wire tmp45;
    wire tmp46;
    wire tmp47;
    wire tmp48;
    wire tmp49;
    wire tmp50;
    wire tmp51;
    wire tmp52;
    wire tmp53;
    wire tmp54;
    wire tmp55;
    wire tmp56;
    wire tmp57;
    wire tmp58;
    wire tmp59;
    wire tmp60;
    wire tmp61;
    wire tmp62;
    wire tmp63;
    wire tmp64;
    wire[63:0] tmp65;
    wire[63:0] tmp66;
    wire tmp67;
    wire tmp68;
    wire[62:0] tmp69;
    wire[63:0] tmp70;
    wire[63:0] tmp71;
    wire tmp72;
    wire tmp73;
    wire tmp74;
    wire tmp75;
    wire tmp76;
    wire tmp77;
    wire[61:0] tmp78;
    wire[63:0] tmp79;
    wire[63:0] tmp80;
    wire tmp81;
    wire tmp82;
    wire[1:0] tmp83;
    wire tmp84;
    wire[1:0] tmp85;
    wire[1:0] tmp86;
    wire tmp87;
    wire tmp88;
    wire[59:0] tmp89;
    wire[63:0] tmp90;
    wire[63:0] tmp91;
    wire tmp92;
    wire tmp93;
    wire[3:0] tmp94;
    wire[2:0] tmp95;
    wire[3:0] tmp96;
    wire[3:0] tmp97;
    wire tmp98;
    wire tmp99;
    wire[55:0] tmp100;
    wire[63:0] tmp101;
    wire[63:0] tmp102;
    wire tmp103;
    wire tmp104;
    wire[7:0] tmp105;
    wire[6:0] tmp106;
    wire[7:0] tmp107;
    wire[7:0] tmp108;
    wire tmp109;
    wire tmp110;
    wire[47:0] tmp111;
    wire[63:0] tmp112;
    wire[63:0] tmp113;
    wire tmp114;
    wire tmp115;
    wire[15:0] tmp116;
    wire[14:0] tmp117;
    wire[15:0] tmp118;
    wire[15:0] tmp119;
    wire tmp120;
    wire tmp121;
    wire[31:0] tmp122;
    wire[63:0] tmp123;
    wire[63:0] tmp124;
    wire tmp125;
    wire tmp126;
    wire[31:0] tmp127;
    wire[30:0] tmp128;
    wire[31:0] tmp129;
    wire[31:0] tmp130;
    wire tmp131;
    wire tmp132;
    wire tmp133;
    wire tmp134;
    wire tmp135;
    wire tmp136;
    wire tmp137;
    wire tmp138;
    wire tmp139;
    wire tmp140;
    wire tmp141;
    wire tmp142;
    wire tmp143;
    wire tmp144;
    wire tmp145;
    wire tmp146;
    wire tmp147;
    wire tmp148;
    wire tmp149;
    wire tmp150;
    wire tmp151;
    wire tmp152;
    wire tmp153;
    wire tmp154;
    wire tmp155;
    wire tmp156;
    wire tmp157;
    wire tmp158;
    wire tmp159;
    wire tmp160;
    wire tmp161;
    wire tmp162;
    wire tmp163;
    wire tmp164;
    wire tmp165;
    wire tmp166;
    wire tmp167;
    wire tmp168;
    wire tmp169;
    wire tmp170;
    wire tmp171;
    wire tmp172;
    wire tmp173;
    wire tmp174;
    wire tmp175;
    wire tmp176;
    wire tmp177;
    wire tmp178;
    wire tmp179;
    wire tmp180;
    wire tmp181;
    wire tmp182;
    wire tmp183;
    wire tmp184;
    wire tmp185;
    wire tmp186;
    wire tmp187;
    wire tmp188;
    wire tmp189;
    wire tmp190;
    wire tmp191;
    wire tmp192;
    wire tmp193;
    wire tmp194;
    wire tmp195;
    wire[63:0] tmp196;
    wire[63:0] tmp197;
    wire[63:0] tmp198;
    wire[63:0] tmp199;
    wire[15:0] tmp200;
    wire[7:0] tmp201;
    wire[3:0] tmp202;
    wire[1:0] tmp203;
    wire tmp204;
    wire tmp205;
    wire tmp206;
    wire tmp207;
    wire tmp208;
    wire[1:0] tmp209;
    wire tmp210;
    wire tmp211;
    wire tmp212;
    wire tmp213;
    wire tmp214;
    wire tmp215;
    wire[3:0] tmp216;
    wire[1:0] tmp217;
    wire tmp218;
    wire tmp219;
    wire tmp220;
    wire tmp221;
    wire tmp222;
    wire[1:0] tmp223;
    wire tmp224;
    wire tmp225;
    wire tmp226;
    wire tmp227;
    wire tmp228;
    wire tmp229;
    wire tmp230;
    wire[7:0] tmp231;
    wire[3:0] tmp232;
    wire[1:0] tmp233;
    wire tmp234;
    wire tmp235;
    wire tmp236;
    wire tmp237;
    wire tmp238;
    wire[1:0] tmp239;
    wire tmp240;
    wire tmp241;
    wire tmp242;
    wire tmp243;
    wire tmp244;
    wire tmp245;
    wire[3:0] tmp246;
    wire[1:0] tmp247;
    wire tmp248;
    wire tmp249;
    wire tmp250;
    wire tmp251;
    wire tmp252;
    wire[1:0] tmp253;
    wire tmp254;
    wire tmp255;
    wire tmp256;
    wire tmp257;
    wire tmp258;
    wire tmp259;
    wire tmp260;
    wire tmp261;
    wire[15:0] tmp262;
    wire[7:0] tmp263;
    wire[3:0] tmp264;
    wire[1:0] tmp265;
    wire tmp266;
    wire tmp267;
    wire tmp268;
    wire tmp269;
    wire tmp270;
    wire[1:0] tmp271;
    wire tmp272;
    wire tmp273;
    wire tmp274;
    wire tmp275;
    wire tmp276;
    wire tmp277;
    wire[3:0] tmp278;
    wire[1:0] tmp279;
    wire tmp280;
    wire tmp281;
    wire tmp282;
    wire tmp283;
    wire tmp284;
    wire[1:0] tmp285;
    wire tmp286;
    wire tmp287;
    wire tmp288;
    wire tmp289;
    wire tmp290;
    wire tmp291;
    wire tmp292;
    wire[7:0] tmp293;
    wire[3:0] tmp294;
    wire[1:0] tmp295;
    wire tmp296;
    wire tmp297;
    wire tmp298;
    wire tmp299;
    wire tmp300;
    wire[1:0] tmp301;
    wire tmp302;
    wire tmp303;
    wire tmp304;
    wire tmp305;
    wire tmp306;
    wire tmp307;
    wire[3:0] tmp308;
    wire[1:0] tmp309;
    wire tmp310;
    wire tmp311;
    wire tmp312;
    wire tmp313;
    wire tmp314;
    wire[1:0] tmp315;
    wire tmp316;
    wire tmp317;
    wire tmp318;
    wire tmp319;
    wire tmp320;
    wire tmp321;
    wire tmp322;
    wire tmp323;
    wire tmp324;
    wire[7:0] tmp325;
    wire[3:0] tmp326;
    wire[1:0] tmp327;
    wire tmp328;
    wire tmp329;
    wire tmp330;
    wire tmp331;
    wire tmp332;
    wire[1:0] tmp333;
    wire tmp334;
    wire tmp335;
    wire tmp336;
    wire tmp337;
    wire tmp338;
    wire tmp339;
    wire[3:0] tmp340;
    wire[1:0] tmp341;
    wire tmp342;
    wire tmp343;
    wire tmp344;
    wire tmp345;
    wire tmp346;
    wire[1:0] tmp347;
    wire tmp348;
    wire tmp349;
    wire tmp350;
    wire tmp351;
    wire tmp352;
    wire tmp353;
    wire tmp354;
    wire[7:0] tmp355;
    wire[3:0] tmp356;
    wire[1:0] tmp357;
    wire tmp358;
    wire tmp359;
    wire tmp360;
    wire tmp361;
    wire tmp362;
    wire[1:0] tmp363;
    wire tmp364;
    wire tmp365;
    wire tmp366;
    wire tmp367;
    wire tmp368;
    wire tmp369;
    wire[3:0] tmp370;
    wire[1:0] tmp371;
    wire tmp372;
    wire tmp373;
    wire tmp374;
    wire tmp375;
    wire tmp376;
    wire[1:0] tmp377;
    wire tmp378;
    wire tmp379;
    wire tmp380;
    wire tmp381;
    wire tmp382;
    wire tmp383;
    wire tmp384;
    wire tmp385;
    wire tmp386;
    wire[3:0] tmp387;
    wire[1:0] tmp388;
    wire tmp389;
    wire tmp390;
    wire tmp391;
    wire tmp392;
    wire tmp393;
    wire[1:0] tmp394;
    wire tmp395;
    wire tmp396;
    wire tmp397;
    wire tmp398;
    wire tmp399;
    wire tmp400;
    wire[3:0] tmp401;
    wire[1:0] tmp402;
    wire tmp403;
    wire tmp404;
    wire tmp405;
    wire tmp406;
    wire tmp407;
    wire[1:0] tmp408;
    wire tmp409;
    wire tmp410;
    wire tmp411;
    wire tmp412;
    wire tmp413;
    wire tmp414;
    wire tmp415;
    wire tmp416;
    wire[1:0] tmp417;
    wire tmp418;
    wire tmp419;
    wire tmp420;
    wire tmp421;
    wire tmp422;
    wire[1:0] tmp423;
    wire tmp424;
    wire tmp425;
    wire tmp426;
    wire tmp427;
    wire tmp428;
    wire tmp429;
    wire tmp430;
    wire tmp431;
    wire tmp432;
    wire tmp433;
    wire tmp434;
    wire tmp435;
    wire tmp436;
    wire tmp437;
    wire tmp438;

    // Combinational
    assign const_0_0 = 0;
    assign const_1_0 = 0;
    assign const_2_0 = 0;
    assign const_3_0 = 0;
    assign const_4_0 = 0;
    assign const_5_0 = 0;
    assign const_6_0 = 0;
    assign const_7_0 = 0;
    assign const_8_0 = 0;
    assign const_9_0 = 0;
    assign const_10_0 = 0;
    assign const_11_0 = 0;
    assign const_12_0 = 0;
    assign const_13_0 = 0;
    assign const_14_0 = 0;
    assign const_15_0 = 0;
    assign const_16_0 = 0;
    assign const_17_0 = 0;
    assign const_18_0 = 0;
    assign const_19_0 = 0;
    assign const_20_0 = 0;
    assign const_21_0 = 0;
    assign const_22_0 = 0;
    assign const_23_0 = 0;
    assign const_24_0 = 0;
    assign overflow = tmp438;
    assign reverse_in = tmp66;
    assign reverse_out = tmp197;
    assign s = tmp199;
    assign shift_1 = tmp71;
    assign shift_2 = tmp80;
    assign shift_4 = tmp91;
    assign shift_8 = tmp102;
    assign shift_16 = tmp113;
    assign shift_32 = tmp124;
    assign shift_off_1 = tmp75;
    assign shift_off_2 = tmp86;
    assign shift_off_4 = tmp97;
    assign shift_off_8 = tmp108;
    assign shift_off_16 = tmp119;
    assign shift_off_32 = tmp130;
    assign tmp0 = direction == const_0_0;
    assign tmp1 = {a[63]};
    assign tmp2 = {a[62]};
    assign tmp3 = {a[61]};
    assign tmp4 = {a[60]};
    assign tmp5 = {a[59]};
    assign tmp6 = {a[58]};
    assign tmp7 = {a[57]};
    assign tmp8 = {a[56]};
    assign tmp9 = {a[55]};
    assign tmp10 = {a[54]};
    assign tmp11 = {a[53]};
    assign tmp12 = {a[52]};
    assign tmp13 = {a[51]};
    assign tmp14 = {a[50]};
    assign tmp15 = {a[49]};
    assign tmp16 = {a[48]};
    assign tmp17 = {a[47]};
    assign tmp18 = {a[46]};
    assign tmp19 = {a[45]};
    assign tmp20 = {a[44]};
    assign tmp21 = {a[43]};
    assign tmp22 = {a[42]};
    assign tmp23 = {a[41]};
    assign tmp24 = {a[40]};
    assign tmp25 = {a[39]};
    assign tmp26 = {a[38]};
    assign tmp27 = {a[37]};
    assign tmp28 = {a[36]};
    assign tmp29 = {a[35]};
    assign tmp30 = {a[34]};
    assign tmp31 = {a[33]};
    assign tmp32 = {a[32]};
    assign tmp33 = {a[31]};
    assign tmp34 = {a[30]};
    assign tmp35 = {a[29]};
    assign tmp36 = {a[28]};
    assign tmp37 = {a[27]};
    assign tmp38 = {a[26]};
    assign tmp39 = {a[25]};
    assign tmp40 = {a[24]};
    assign tmp41 = {a[23]};
    assign tmp42 = {a[22]};
    assign tmp43 = {a[21]};
    assign tmp44 = {a[20]};
    assign tmp45 = {a[19]};
    assign tmp46 = {a[18]};
    assign tmp47 = {a[17]};
    assign tmp48 = {a[16]};
    assign tmp49 = {a[15]};
    assign tmp50 = {a[14]};
    assign tmp51 = {a[13]};
    assign tmp52 = {a[12]};
    assign tmp53 = {a[11]};
    assign tmp54 = {a[10]};
    assign tmp55 = {a[9]};
    assign tmp56 = {a[8]};
    assign tmp57 = {a[7]};
    assign tmp58 = {a[6]};
    assign tmp59 = {a[5]};
    assign tmp60 = {a[4]};
    assign tmp61 = {a[3]};
    assign tmp62 = {a[2]};
    assign tmp63 = {a[1]};
    assign tmp64 = {a[0]};
    assign tmp65 = {tmp64, tmp63, tmp62, tmp61, tmp60, tmp59, tmp58, tmp57, tmp56, tmp55, tmp54, tmp53, tmp52, tmp51, tmp50, tmp49, tmp48, tmp47, tmp46, tmp45, tmp44, tmp43, tmp42, tmp41, tmp40, tmp39, tmp38, tmp37, tmp36, tmp35, tmp34, tmp33, tmp32, tmp31, tmp30, tmp29, tmp28, tmp27, tmp26, tmp25, tmp24, tmp23, tmp22, tmp21, tmp20, tmp19, tmp18, tmp17, tmp16, tmp15, tmp14, tmp13, tmp12, tmp11, tmp10, tmp9, tmp8, tmp7, tmp6, tmp5, tmp4, tmp3, tmp2, tmp1};
    assign tmp66 = tmp0 ? a : tmp65;
    assign tmp67 = {n[0]};
    assign tmp68 = tmp67 == const_1_0;
    assign tmp69 = {reverse_in[62], reverse_in[61], reverse_in[60], reverse_in[59], reverse_in[58], reverse_in[57], reverse_in[56], reverse_in[55], reverse_in[54], reverse_in[53], reverse_in[52], reverse_in[51], reverse_in[50], reverse_in[49], reverse_in[48], reverse_in[47], reverse_in[46], reverse_in[45], reverse_in[44], reverse_in[43], reverse_in[42], reverse_in[41], reverse_in[40], reverse_in[39], reverse_in[38], reverse_in[37], reverse_in[36], reverse_in[35], reverse_in[34], reverse_in[33], reverse_in[32], reverse_in[31], reverse_in[30], reverse_in[29], reverse_in[28], reverse_in[27], reverse_in[26], reverse_in[25], reverse_in[24], reverse_in[23], reverse_in[22], reverse_in[21], reverse_in[20], reverse_in[19], reverse_in[18], reverse_in[17], reverse_in[16], reverse_in[15], reverse_in[14], reverse_in[13], reverse_in[12], reverse_in[11], reverse_in[10], reverse_in[9], reverse_in[8], reverse_in[7], reverse_in[6], reverse_in[5], reverse_in[4], reverse_in[3], reverse_in[2], reverse_in[1], reverse_in[0]};
    assign tmp70 = {tmp69, shift_in};
    assign tmp71 = tmp68 ? reverse_in : tmp70;
    assign tmp72 = {n[0]};
    assign tmp73 = tmp72 == const_2_0;
    assign tmp74 = {reverse_in[63]};
    assign tmp75 = tmp73 ? const_3_0 : tmp74;
    assign tmp76 = {n[1]};
    assign tmp77 = tmp76 == const_4_0;
    assign tmp78 = {shift_1[61], shift_1[60], shift_1[59], shift_1[58], shift_1[57], shift_1[56], shift_1[55], shift_1[54], shift_1[53], shift_1[52], shift_1[51], shift_1[50], shift_1[49], shift_1[48], shift_1[47], shift_1[46], shift_1[45], shift_1[44], shift_1[43], shift_1[42], shift_1[41], shift_1[40], shift_1[39], shift_1[38], shift_1[37], shift_1[36], shift_1[35], shift_1[34], shift_1[33], shift_1[32], shift_1[31], shift_1[30], shift_1[29], shift_1[28], shift_1[27], shift_1[26], shift_1[25], shift_1[24], shift_1[23], shift_1[22], shift_1[21], shift_1[20], shift_1[19], shift_1[18], shift_1[17], shift_1[16], shift_1[15], shift_1[14], shift_1[13], shift_1[12], shift_1[11], shift_1[10], shift_1[9], shift_1[8], shift_1[7], shift_1[6], shift_1[5], shift_1[4], shift_1[3], shift_1[2], shift_1[1], shift_1[0]};
    assign tmp79 = {tmp78, shift_in, shift_in};
    assign tmp80 = tmp77 ? shift_1 : tmp79;
    assign tmp81 = {n[1]};
    assign tmp82 = tmp81 == const_5_0;
    assign tmp83 = {shift_1[63], shift_1[62]};
    assign tmp84 = {const_7_0};
    assign tmp85 = {tmp84, const_6_0};
    assign tmp86 = tmp82 ? tmp85 : tmp83;
    assign tmp87 = {n[2]};
    assign tmp88 = tmp87 == const_8_0;
    assign tmp89 = {shift_2[59], shift_2[58], shift_2[57], shift_2[56], shift_2[55], shift_2[54], shift_2[53], shift_2[52], shift_2[51], shift_2[50], shift_2[49], shift_2[48], shift_2[47], shift_2[46], shift_2[45], shift_2[44], shift_2[43], shift_2[42], shift_2[41], shift_2[40], shift_2[39], shift_2[38], shift_2[37], shift_2[36], shift_2[35], shift_2[34], shift_2[33], shift_2[32], shift_2[31], shift_2[30], shift_2[29], shift_2[28], shift_2[27], shift_2[26], shift_2[25], shift_2[24], shift_2[23], shift_2[22], shift_2[21], shift_2[20], shift_2[19], shift_2[18], shift_2[17], shift_2[16], shift_2[15], shift_2[14], shift_2[13], shift_2[12], shift_2[11], shift_2[10], shift_2[9], shift_2[8], shift_2[7], shift_2[6], shift_2[5], shift_2[4], shift_2[3], shift_2[2], shift_2[1], shift_2[0]};
    assign tmp90 = {tmp89, shift_in, shift_in, shift_in, shift_in};
    assign tmp91 = tmp88 ? shift_2 : tmp90;
    assign tmp92 = {n[1]};
    assign tmp93 = tmp92 == const_9_0;
    assign tmp94 = {shift_2[63], shift_2[62], shift_2[61], shift_2[60]};
    assign tmp95 = {const_11_0, const_11_0, const_11_0};
    assign tmp96 = {tmp95, const_10_0};
    assign tmp97 = tmp93 ? tmp96 : tmp94;
    assign tmp98 = {n[3]};
    assign tmp99 = tmp98 == const_12_0;
    assign tmp100 = {shift_4[55], shift_4[54], shift_4[53], shift_4[52], shift_4[51], shift_4[50], shift_4[49], shift_4[48], shift_4[47], shift_4[46], shift_4[45], shift_4[44], shift_4[43], shift_4[42], shift_4[41], shift_4[40], shift_4[39], shift_4[38], shift_4[37], shift_4[36], shift_4[35], shift_4[34], shift_4[33], shift_4[32], shift_4[31], shift_4[30], shift_4[29], shift_4[28], shift_4[27], shift_4[26], shift_4[25], shift_4[24], shift_4[23], shift_4[22], shift_4[21], shift_4[20], shift_4[19], shift_4[18], shift_4[17], shift_4[16], shift_4[15], shift_4[14], shift_4[13], shift_4[12], shift_4[11], shift_4[10], shift_4[9], shift_4[8], shift_4[7], shift_4[6], shift_4[5], shift_4[4], shift_4[3], shift_4[2], shift_4[1], shift_4[0]};
    assign tmp101 = {tmp100, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in};
    assign tmp102 = tmp99 ? shift_4 : tmp101;
    assign tmp103 = {n[1]};
    assign tmp104 = tmp103 == const_13_0;
    assign tmp105 = {shift_4[63], shift_4[62], shift_4[61], shift_4[60], shift_4[59], shift_4[58], shift_4[57], shift_4[56]};
    assign tmp106 = {const_15_0, const_15_0, const_15_0, const_15_0, const_15_0, const_15_0, const_15_0};
    assign tmp107 = {tmp106, const_14_0};
    assign tmp108 = tmp104 ? tmp107 : tmp105;
    assign tmp109 = {n[4]};
    assign tmp110 = tmp109 == const_16_0;
    assign tmp111 = {shift_8[47], shift_8[46], shift_8[45], shift_8[44], shift_8[43], shift_8[42], shift_8[41], shift_8[40], shift_8[39], shift_8[38], shift_8[37], shift_8[36], shift_8[35], shift_8[34], shift_8[33], shift_8[32], shift_8[31], shift_8[30], shift_8[29], shift_8[28], shift_8[27], shift_8[26], shift_8[25], shift_8[24], shift_8[23], shift_8[22], shift_8[21], shift_8[20], shift_8[19], shift_8[18], shift_8[17], shift_8[16], shift_8[15], shift_8[14], shift_8[13], shift_8[12], shift_8[11], shift_8[10], shift_8[9], shift_8[8], shift_8[7], shift_8[6], shift_8[5], shift_8[4], shift_8[3], shift_8[2], shift_8[1], shift_8[0]};
    assign tmp112 = {tmp111, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in};
    assign tmp113 = tmp110 ? shift_8 : tmp112;
    assign tmp114 = {n[1]};
    assign tmp115 = tmp114 == const_17_0;
    assign tmp116 = {shift_8[63], shift_8[62], shift_8[61], shift_8[60], shift_8[59], shift_8[58], shift_8[57], shift_8[56], shift_8[55], shift_8[54], shift_8[53], shift_8[52], shift_8[51], shift_8[50], shift_8[49], shift_8[48]};
    assign tmp117 = {const_19_0, const_19_0, const_19_0, const_19_0, const_19_0, const_19_0, const_19_0, const_19_0, const_19_0, const_19_0, const_19_0, const_19_0, const_19_0, const_19_0, const_19_0};
    assign tmp118 = {tmp117, const_18_0};
    assign tmp119 = tmp115 ? tmp118 : tmp116;
    assign tmp120 = {n[5]};
    assign tmp121 = tmp120 == const_20_0;
    assign tmp122 = {shift_16[31], shift_16[30], shift_16[29], shift_16[28], shift_16[27], shift_16[26], shift_16[25], shift_16[24], shift_16[23], shift_16[22], shift_16[21], shift_16[20], shift_16[19], shift_16[18], shift_16[17], shift_16[16], shift_16[15], shift_16[14], shift_16[13], shift_16[12], shift_16[11], shift_16[10], shift_16[9], shift_16[8], shift_16[7], shift_16[6], shift_16[5], shift_16[4], shift_16[3], shift_16[2], shift_16[1], shift_16[0]};
    assign tmp123 = {tmp122, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in};
    assign tmp124 = tmp121 ? shift_16 : tmp123;
    assign tmp125 = {n[1]};
    assign tmp126 = tmp125 == const_21_0;
    assign tmp127 = {shift_16[63], shift_16[62], shift_16[61], shift_16[60], shift_16[59], shift_16[58], shift_16[57], shift_16[56], shift_16[55], shift_16[54], shift_16[53], shift_16[52], shift_16[51], shift_16[50], shift_16[49], shift_16[48], shift_16[47], shift_16[46], shift_16[45], shift_16[44], shift_16[43], shift_16[42], shift_16[41], shift_16[40], shift_16[39], shift_16[38], shift_16[37], shift_16[36], shift_16[35], shift_16[34], shift_16[33], shift_16[32]};
    assign tmp128 = {const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0};
    assign tmp129 = {tmp128, const_22_0};
    assign tmp130 = tmp126 ? tmp129 : tmp127;
    assign tmp131 = direction == const_24_0;
    assign tmp132 = {shift_32[63]};
    assign tmp133 = {shift_32[62]};
    assign tmp134 = {shift_32[61]};
    assign tmp135 = {shift_32[60]};
    assign tmp136 = {shift_32[59]};
    assign tmp137 = {shift_32[58]};
    assign tmp138 = {shift_32[57]};
    assign tmp139 = {shift_32[56]};
    assign tmp140 = {shift_32[55]};
    assign tmp141 = {shift_32[54]};
    assign tmp142 = {shift_32[53]};
    assign tmp143 = {shift_32[52]};
    assign tmp144 = {shift_32[51]};
    assign tmp145 = {shift_32[50]};
    assign tmp146 = {shift_32[49]};
    assign tmp147 = {shift_32[48]};
    assign tmp148 = {shift_32[47]};
    assign tmp149 = {shift_32[46]};
    assign tmp150 = {shift_32[45]};
    assign tmp151 = {shift_32[44]};
    assign tmp152 = {shift_32[43]};
    assign tmp153 = {shift_32[42]};
    assign tmp154 = {shift_32[41]};
    assign tmp155 = {shift_32[40]};
    assign tmp156 = {shift_32[39]};
    assign tmp157 = {shift_32[38]};
    assign tmp158 = {shift_32[37]};
    assign tmp159 = {shift_32[36]};
    assign tmp160 = {shift_32[35]};
    assign tmp161 = {shift_32[34]};
    assign tmp162 = {shift_32[33]};
    assign tmp163 = {shift_32[32]};
    assign tmp164 = {shift_32[31]};
    assign tmp165 = {shift_32[30]};
    assign tmp166 = {shift_32[29]};
    assign tmp167 = {shift_32[28]};
    assign tmp168 = {shift_32[27]};
    assign tmp169 = {shift_32[26]};
    assign tmp170 = {shift_32[25]};
    assign tmp171 = {shift_32[24]};
    assign tmp172 = {shift_32[23]};
    assign tmp173 = {shift_32[22]};
    assign tmp174 = {shift_32[21]};
    assign tmp175 = {shift_32[20]};
    assign tmp176 = {shift_32[19]};
    assign tmp177 = {shift_32[18]};
    assign tmp178 = {shift_32[17]};
    assign tmp179 = {shift_32[16]};
    assign tmp180 = {shift_32[15]};
    assign tmp181 = {shift_32[14]};
    assign tmp182 = {shift_32[13]};
    assign tmp183 = {shift_32[12]};
    assign tmp184 = {shift_32[11]};
    assign tmp185 = {shift_32[10]};
    assign tmp186 = {shift_32[9]};
    assign tmp187 = {shift_32[8]};
    assign tmp188 = {shift_32[7]};
    assign tmp189 = {shift_32[6]};
    assign tmp190 = {shift_32[5]};
    assign tmp191 = {shift_32[4]};
    assign tmp192 = {shift_32[3]};
    assign tmp193 = {shift_32[2]};
    assign tmp194 = {shift_32[1]};
    assign tmp195 = {shift_32[0]};
    assign tmp196 = {tmp195, tmp194, tmp193, tmp192, tmp191, tmp190, tmp189, tmp188, tmp187, tmp186, tmp185, tmp184, tmp183, tmp182, tmp181, tmp180, tmp179, tmp178, tmp177, tmp176, tmp175, tmp174, tmp173, tmp172, tmp171, tmp170, tmp169, tmp168, tmp167, tmp166, tmp165, tmp164, tmp163, tmp162, tmp161, tmp160, tmp159, tmp158, tmp157, tmp156, tmp155, tmp154, tmp153, tmp152, tmp151, tmp150, tmp149, tmp148, tmp147, tmp146, tmp145, tmp144, tmp143, tmp142, tmp141, tmp140, tmp139, tmp138, tmp137, tmp136, tmp135, tmp134, tmp133, tmp132};
    assign tmp197 = tmp131 ? shift_32 : tmp196;
    assign tmp198 = ~reverse_out;
    assign tmp199 = invert ? tmp198 : reverse_out;
    assign tmp200 = {shift_off_32[15], shift_off_32[14], shift_off_32[13], shift_off_32[12], shift_off_32[11], shift_off_32[10], shift_off_32[9], shift_off_32[8], shift_off_32[7], shift_off_32[6], shift_off_32[5], shift_off_32[4], shift_off_32[3], shift_off_32[2], shift_off_32[1], shift_off_32[0]};
    assign tmp201 = {tmp200[7], tmp200[6], tmp200[5], tmp200[4], tmp200[3], tmp200[2], tmp200[1], tmp200[0]};
    assign tmp202 = {tmp201[3], tmp201[2], tmp201[1], tmp201[0]};
    assign tmp203 = {tmp202[1], tmp202[0]};
    assign tmp204 = {tmp203[0]};
    assign tmp205 = {tmp204};
    assign tmp206 = {tmp203[1]};
    assign tmp207 = {tmp206};
    assign tmp208 = tmp205 | tmp207;
    assign tmp209 = {tmp202[3], tmp202[2]};
    assign tmp210 = {tmp209[0]};
    assign tmp211 = {tmp210};
    assign tmp212 = {tmp209[1]};
    assign tmp213 = {tmp212};
    assign tmp214 = tmp211 | tmp213;
    assign tmp215 = tmp208 | tmp214;
    assign tmp216 = {tmp201[7], tmp201[6], tmp201[5], tmp201[4]};
    assign tmp217 = {tmp216[1], tmp216[0]};
    assign tmp218 = {tmp217[0]};
    assign tmp219 = {tmp218};
    assign tmp220 = {tmp217[1]};
    assign tmp221 = {tmp220};
    assign tmp222 = tmp219 | tmp221;
    assign tmp223 = {tmp216[3], tmp216[2]};
    assign tmp224 = {tmp223[0]};
    assign tmp225 = {tmp224};
    assign tmp226 = {tmp223[1]};
    assign tmp227 = {tmp226};
    assign tmp228 = tmp225 | tmp227;
    assign tmp229 = tmp222 | tmp228;
    assign tmp230 = tmp215 | tmp229;
    assign tmp231 = {tmp200[15], tmp200[14], tmp200[13], tmp200[12], tmp200[11], tmp200[10], tmp200[9], tmp200[8]};
    assign tmp232 = {tmp231[3], tmp231[2], tmp231[1], tmp231[0]};
    assign tmp233 = {tmp232[1], tmp232[0]};
    assign tmp234 = {tmp233[0]};
    assign tmp235 = {tmp234};
    assign tmp236 = {tmp233[1]};
    assign tmp237 = {tmp236};
    assign tmp238 = tmp235 | tmp237;
    assign tmp239 = {tmp232[3], tmp232[2]};
    assign tmp240 = {tmp239[0]};
    assign tmp241 = {tmp240};
    assign tmp242 = {tmp239[1]};
    assign tmp243 = {tmp242};
    assign tmp244 = tmp241 | tmp243;
    assign tmp245 = tmp238 | tmp244;
    assign tmp246 = {tmp231[7], tmp231[6], tmp231[5], tmp231[4]};
    assign tmp247 = {tmp246[1], tmp246[0]};
    assign tmp248 = {tmp247[0]};
    assign tmp249 = {tmp248};
    assign tmp250 = {tmp247[1]};
    assign tmp251 = {tmp250};
    assign tmp252 = tmp249 | tmp251;
    assign tmp253 = {tmp246[3], tmp246[2]};
    assign tmp254 = {tmp253[0]};
    assign tmp255 = {tmp254};
    assign tmp256 = {tmp253[1]};
    assign tmp257 = {tmp256};
    assign tmp258 = tmp255 | tmp257;
    assign tmp259 = tmp252 | tmp258;
    assign tmp260 = tmp245 | tmp259;
    assign tmp261 = tmp230 | tmp260;
    assign tmp262 = {shift_off_32[31], shift_off_32[30], shift_off_32[29], shift_off_32[28], shift_off_32[27], shift_off_32[26], shift_off_32[25], shift_off_32[24], shift_off_32[23], shift_off_32[22], shift_off_32[21], shift_off_32[20], shift_off_32[19], shift_off_32[18], shift_off_32[17], shift_off_32[16]};
    assign tmp263 = {tmp262[7], tmp262[6], tmp262[5], tmp262[4], tmp262[3], tmp262[2], tmp262[1], tmp262[0]};
    assign tmp264 = {tmp263[3], tmp263[2], tmp263[1], tmp263[0]};
    assign tmp265 = {tmp264[1], tmp264[0]};
    assign tmp266 = {tmp265[0]};
    assign tmp267 = {tmp266};
    assign tmp268 = {tmp265[1]};
    assign tmp269 = {tmp268};
    assign tmp270 = tmp267 | tmp269;
    assign tmp271 = {tmp264[3], tmp264[2]};
    assign tmp272 = {tmp271[0]};
    assign tmp273 = {tmp272};
    assign tmp274 = {tmp271[1]};
    assign tmp275 = {tmp274};
    assign tmp276 = tmp273 | tmp275;
    assign tmp277 = tmp270 | tmp276;
    assign tmp278 = {tmp263[7], tmp263[6], tmp263[5], tmp263[4]};
    assign tmp279 = {tmp278[1], tmp278[0]};
    assign tmp280 = {tmp279[0]};
    assign tmp281 = {tmp280};
    assign tmp282 = {tmp279[1]};
    assign tmp283 = {tmp282};
    assign tmp284 = tmp281 | tmp283;
    assign tmp285 = {tmp278[3], tmp278[2]};
    assign tmp286 = {tmp285[0]};
    assign tmp287 = {tmp286};
    assign tmp288 = {tmp285[1]};
    assign tmp289 = {tmp288};
    assign tmp290 = tmp287 | tmp289;
    assign tmp291 = tmp284 | tmp290;
    assign tmp292 = tmp277 | tmp291;
    assign tmp293 = {tmp262[15], tmp262[14], tmp262[13], tmp262[12], tmp262[11], tmp262[10], tmp262[9], tmp262[8]};
    assign tmp294 = {tmp293[3], tmp293[2], tmp293[1], tmp293[0]};
    assign tmp295 = {tmp294[1], tmp294[0]};
    assign tmp296 = {tmp295[0]};
    assign tmp297 = {tmp296};
    assign tmp298 = {tmp295[1]};
    assign tmp299 = {tmp298};
    assign tmp300 = tmp297 | tmp299;
    assign tmp301 = {tmp294[3], tmp294[2]};
    assign tmp302 = {tmp301[0]};
    assign tmp303 = {tmp302};
    assign tmp304 = {tmp301[1]};
    assign tmp305 = {tmp304};
    assign tmp306 = tmp303 | tmp305;
    assign tmp307 = tmp300 | tmp306;
    assign tmp308 = {tmp293[7], tmp293[6], tmp293[5], tmp293[4]};
    assign tmp309 = {tmp308[1], tmp308[0]};
    assign tmp310 = {tmp309[0]};
    assign tmp311 = {tmp310};
    assign tmp312 = {tmp309[1]};
    assign tmp313 = {tmp312};
    assign tmp314 = tmp311 | tmp313;
    assign tmp315 = {tmp308[3], tmp308[2]};
    assign tmp316 = {tmp315[0]};
    assign tmp317 = {tmp316};
    assign tmp318 = {tmp315[1]};
    assign tmp319 = {tmp318};
    assign tmp320 = tmp317 | tmp319;
    assign tmp321 = tmp314 | tmp320;
    assign tmp322 = tmp307 | tmp321;
    assign tmp323 = tmp292 | tmp322;
    assign tmp324 = tmp261 | tmp323;
    assign tmp325 = {shift_off_16[7], shift_off_16[6], shift_off_16[5], shift_off_16[4], shift_off_16[3], shift_off_16[2], shift_off_16[1], shift_off_16[0]};
    assign tmp326 = {tmp325[3], tmp325[2], tmp325[1], tmp325[0]};
    assign tmp327 = {tmp326[1], tmp326[0]};
    assign tmp328 = {tmp327[0]};
    assign tmp329 = {tmp328};
    assign tmp330 = {tmp327[1]};
    assign tmp331 = {tmp330};
    assign tmp332 = tmp329 | tmp331;
    assign tmp333 = {tmp326[3], tmp326[2]};
    assign tmp334 = {tmp333[0]};
    assign tmp335 = {tmp334};
    assign tmp336 = {tmp333[1]};
    assign tmp337 = {tmp336};
    assign tmp338 = tmp335 | tmp337;
    assign tmp339 = tmp332 | tmp338;
    assign tmp340 = {tmp325[7], tmp325[6], tmp325[5], tmp325[4]};
    assign tmp341 = {tmp340[1], tmp340[0]};
    assign tmp342 = {tmp341[0]};
    assign tmp343 = {tmp342};
    assign tmp344 = {tmp341[1]};
    assign tmp345 = {tmp344};
    assign tmp346 = tmp343 | tmp345;
    assign tmp347 = {tmp340[3], tmp340[2]};
    assign tmp348 = {tmp347[0]};
    assign tmp349 = {tmp348};
    assign tmp350 = {tmp347[1]};
    assign tmp351 = {tmp350};
    assign tmp352 = tmp349 | tmp351;
    assign tmp353 = tmp346 | tmp352;
    assign tmp354 = tmp339 | tmp353;
    assign tmp355 = {shift_off_16[15], shift_off_16[14], shift_off_16[13], shift_off_16[12], shift_off_16[11], shift_off_16[10], shift_off_16[9], shift_off_16[8]};
    assign tmp356 = {tmp355[3], tmp355[2], tmp355[1], tmp355[0]};
    assign tmp357 = {tmp356[1], tmp356[0]};
    assign tmp358 = {tmp357[0]};
    assign tmp359 = {tmp358};
    assign tmp360 = {tmp357[1]};
    assign tmp361 = {tmp360};
    assign tmp362 = tmp359 | tmp361;
    assign tmp363 = {tmp356[3], tmp356[2]};
    assign tmp364 = {tmp363[0]};
    assign tmp365 = {tmp364};
    assign tmp366 = {tmp363[1]};
    assign tmp367 = {tmp366};
    assign tmp368 = tmp365 | tmp367;
    assign tmp369 = tmp362 | tmp368;
    assign tmp370 = {tmp355[7], tmp355[6], tmp355[5], tmp355[4]};
    assign tmp371 = {tmp370[1], tmp370[0]};
    assign tmp372 = {tmp371[0]};
    assign tmp373 = {tmp372};
    assign tmp374 = {tmp371[1]};
    assign tmp375 = {tmp374};
    assign tmp376 = tmp373 | tmp375;
    assign tmp377 = {tmp370[3], tmp370[2]};
    assign tmp378 = {tmp377[0]};
    assign tmp379 = {tmp378};
    assign tmp380 = {tmp377[1]};
    assign tmp381 = {tmp380};
    assign tmp382 = tmp379 | tmp381;
    assign tmp383 = tmp376 | tmp382;
    assign tmp384 = tmp369 | tmp383;
    assign tmp385 = tmp354 | tmp384;
    assign tmp386 = tmp324 | tmp385;
    assign tmp387 = {shift_off_8[3], shift_off_8[2], shift_off_8[1], shift_off_8[0]};
    assign tmp388 = {tmp387[1], tmp387[0]};
    assign tmp389 = {tmp388[0]};
    assign tmp390 = {tmp389};
    assign tmp391 = {tmp388[1]};
    assign tmp392 = {tmp391};
    assign tmp393 = tmp390 | tmp392;
    assign tmp394 = {tmp387[3], tmp387[2]};
    assign tmp395 = {tmp394[0]};
    assign tmp396 = {tmp395};
    assign tmp397 = {tmp394[1]};
    assign tmp398 = {tmp397};
    assign tmp399 = tmp396 | tmp398;
    assign tmp400 = tmp393 | tmp399;
    assign tmp401 = {shift_off_8[7], shift_off_8[6], shift_off_8[5], shift_off_8[4]};
    assign tmp402 = {tmp401[1], tmp401[0]};
    assign tmp403 = {tmp402[0]};
    assign tmp404 = {tmp403};
    assign tmp405 = {tmp402[1]};
    assign tmp406 = {tmp405};
    assign tmp407 = tmp404 | tmp406;
    assign tmp408 = {tmp401[3], tmp401[2]};
    assign tmp409 = {tmp408[0]};
    assign tmp410 = {tmp409};
    assign tmp411 = {tmp408[1]};
    assign tmp412 = {tmp411};
    assign tmp413 = tmp410 | tmp412;
    assign tmp414 = tmp407 | tmp413;
    assign tmp415 = tmp400 | tmp414;
    assign tmp416 = tmp386 | tmp415;
    assign tmp417 = {shift_off_4[1], shift_off_4[0]};
    assign tmp418 = {tmp417[0]};
    assign tmp419 = {tmp418};
    assign tmp420 = {tmp417[1]};
    assign tmp421 = {tmp420};
    assign tmp422 = tmp419 | tmp421;
    assign tmp423 = {shift_off_4[3], shift_off_4[2]};
    assign tmp424 = {tmp423[0]};
    assign tmp425 = {tmp424};
    assign tmp426 = {tmp423[1]};
    assign tmp427 = {tmp426};
    assign tmp428 = tmp425 | tmp427;
    assign tmp429 = tmp422 | tmp428;
    assign tmp430 = tmp416 | tmp429;
    assign tmp431 = {shift_off_2[0]};
    assign tmp432 = {tmp431};
    assign tmp433 = {shift_off_2[1]};
    assign tmp434 = {tmp433};
    assign tmp435 = tmp432 | tmp434;
    assign tmp436 = tmp430 | tmp435;
    assign tmp437 = {shift_off_1};
    assign tmp438 = tmp436 | tmp437;

endmodule

