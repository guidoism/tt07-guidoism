/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_guidoism (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // All output pins must be assigned. If not used, assign to 0.
  //assign uo_out  = ui_in + uio_in;  // Example: ou_out is the sum of ui_in and uio_in
  //assign uio_out = 0;
  //assign uio_oe  = 0;

// Generated automatically via PyRTL
// As one initial test of synthesis, map to FPGA with:
//   yosys -p "synth_xilinx -top toplevel" thisfile.v
//
// module toplevel(clk, rst, a, direction, invert, n, shift_in, overflow, s);
//    input clk;
//    input rst;
//   
//    input[63:0] a;
//    input direction;
//    input invert;
//    input[5:0] n;
//    input shift_in;
//    output overflow;
//    output[63:0] s;

   wire [63:0]        a;
   assign a[7:0] = ui_in;
   
   wire [5:0]        n;
   wire              direction;
   wire              invert;
   wire              shift_in;
   assign uio_oe = 0;
   assign n[4:0] = uio_in[4:0];
   assign n[5] = 0;
   assign direction = uio_in[5];
   assign invert = uio_in[6];
   assign shift_in = uio_in[7];
   
   wire overflow;
   wire [63:0] s;
   assign s[7:0] = uo_out;
   
    wire const_0_0;
    wire const_1_0;
    wire const_2_0;
    wire const_3_0;
    wire const_4_0;
    wire const_5_0;
    wire const_6_0;
    wire const_7_0;
    wire const_8_0;
    wire const_9_0;
    wire const_10_0;
    wire const_11_0;
    wire const_12_0;
    wire const_13_0;
    wire const_14_0;
    wire const_15_0;
    wire const_16_0;
    wire const_17_0;
    wire const_18_0;
    wire const_19_0;
    wire const_20_0;
    wire const_21_0;
    wire const_22_0;
    wire const_23_0;
    wire const_24_0;
    wire[63:0] reverse_in;
    wire[63:0] reverse_out;
    wire[63:0] shift_1;
    wire[63:0] shift_2;
    wire[63:0] shift_4;
    wire[63:0] shift_8;
    wire[63:0] shift_16;
    wire[63:0] shift_32;
    wire shift_off_1;
    wire[1:0] shift_off_2;
    wire[3:0] shift_off_4;
    wire[7:0] shift_off_8;
    wire[15:0] shift_off_16;
    wire[31:0] shift_off_32;
    wire tmp0_barrel_shifter_line25;
    wire tmp1_barrel_shifter_line25;
    wire tmp2_barrel_shifter_line25;
    wire tmp3_barrel_shifter_line25;
    wire tmp4_barrel_shifter_line25;
    wire tmp5_barrel_shifter_line25;
    wire tmp6_barrel_shifter_line25;
    wire tmp7_barrel_shifter_line25;
    wire tmp8_barrel_shifter_line25;
    wire tmp9_barrel_shifter_line25;
    wire tmp10_barrel_shifter_line25;
    wire tmp11_barrel_shifter_line25;
    wire tmp12_barrel_shifter_line25;
    wire tmp13_barrel_shifter_line25;
    wire tmp14_barrel_shifter_line25;
    wire tmp15_barrel_shifter_line25;
    wire tmp16_barrel_shifter_line25;
    wire tmp17_barrel_shifter_line25;
    wire tmp18_barrel_shifter_line25;
    wire tmp19_barrel_shifter_line25;
    wire tmp20_barrel_shifter_line25;
    wire tmp21_barrel_shifter_line25;
    wire tmp22_barrel_shifter_line25;
    wire tmp23_barrel_shifter_line25;
    wire tmp24_barrel_shifter_line25;
    wire tmp25_barrel_shifter_line25;
    wire tmp26_barrel_shifter_line25;
    wire tmp27_barrel_shifter_line25;
    wire tmp28_barrel_shifter_line25;
    wire tmp29_barrel_shifter_line25;
    wire tmp30_barrel_shifter_line25;
    wire tmp31_barrel_shifter_line25;
    wire tmp32_barrel_shifter_line25;
    wire tmp33_barrel_shifter_line25;
    wire tmp34_barrel_shifter_line25;
    wire tmp35_barrel_shifter_line25;
    wire tmp36_barrel_shifter_line25;
    wire tmp37_barrel_shifter_line25;
    wire tmp38_barrel_shifter_line25;
    wire tmp39_barrel_shifter_line25;
    wire tmp40_barrel_shifter_line25;
    wire tmp41_barrel_shifter_line25;
    wire tmp42_barrel_shifter_line25;
    wire tmp43_barrel_shifter_line25;
    wire tmp44_barrel_shifter_line25;
    wire tmp45_barrel_shifter_line25;
    wire tmp46_barrel_shifter_line25;
    wire tmp47_barrel_shifter_line25;
    wire tmp48_barrel_shifter_line25;
    wire tmp49_barrel_shifter_line25;
    wire tmp50_barrel_shifter_line25;
    wire tmp51_barrel_shifter_line25;
    wire tmp52_barrel_shifter_line25;
    wire tmp53_barrel_shifter_line25;
    wire tmp54_barrel_shifter_line25;
    wire tmp55_barrel_shifter_line25;
    wire tmp56_barrel_shifter_line25;
    wire tmp57_barrel_shifter_line25;
    wire tmp58_barrel_shifter_line25;
    wire tmp59_barrel_shifter_line25;
    wire tmp60_barrel_shifter_line25;
    wire tmp61_barrel_shifter_line25;
    wire tmp62_barrel_shifter_line25;
    wire tmp63_barrel_shifter_line25;
    wire tmp64_barrel_shifter_line25;
    wire[63:0] tmp65_barrel_shifter_line25;
    wire[63:0] tmp66_barrel_shifter_line25;
    wire tmp67_barrel_shifter_line37;
    wire tmp68_barrel_shifter_line37;
    wire[62:0] tmp69_barrel_shifter_line37;
    wire[63:0] tmp70_barrel_shifter_line37;
    wire[63:0] tmp71_barrel_shifter_line37;
    wire tmp72_barrel_shifter_line39;
    wire tmp73_barrel_shifter_line39;
    wire tmp74_barrel_shifter_line39;
    wire tmp75_barrel_shifter_line39;
    wire tmp76_barrel_shifter_line42;
    wire tmp77_barrel_shifter_line42;
    wire[61:0] tmp78_barrel_shifter_line42;
    wire[63:0] tmp79_barrel_shifter_line42;
    wire[63:0] tmp80_barrel_shifter_line42;
    wire tmp81_barrel_shifter_line44;
    wire tmp82_barrel_shifter_line44;
    wire[1:0] tmp83_barrel_shifter_line44;
    wire tmp84_barrel_shifter_line44;
    wire[1:0] tmp85_barrel_shifter_line44;
    wire[1:0] tmp86_barrel_shifter_line44;
    wire tmp87_barrel_shifter_line47;
    wire tmp88_barrel_shifter_line47;
    wire[59:0] tmp89_barrel_shifter_line47;
    wire[63:0] tmp90_barrel_shifter_line47;
    wire[63:0] tmp91_barrel_shifter_line47;
    wire tmp92_barrel_shifter_line49;
    wire tmp93_barrel_shifter_line49;
    wire[3:0] tmp94_barrel_shifter_line49;
    wire[2:0] tmp95_barrel_shifter_line49;
    wire[3:0] tmp96_barrel_shifter_line49;
    wire[3:0] tmp97_barrel_shifter_line49;
    wire tmp98_barrel_shifter_line52;
    wire tmp99_barrel_shifter_line52;
    wire[55:0] tmp100_barrel_shifter_line52;
    wire[63:0] tmp101_barrel_shifter_line52;
    wire[63:0] tmp102_barrel_shifter_line52;
    wire tmp103_barrel_shifter_line54;
    wire tmp104_barrel_shifter_line54;
    wire[7:0] tmp105_barrel_shifter_line54;
    wire[6:0] tmp106_barrel_shifter_line54;
    wire[7:0] tmp107_barrel_shifter_line54;
    wire[7:0] tmp108_barrel_shifter_line54;
    wire tmp109_barrel_shifter_line57;
    wire tmp110_barrel_shifter_line57;
    wire[47:0] tmp111_barrel_shifter_line57;
    wire[63:0] tmp112_barrel_shifter_line57;
    wire[63:0] tmp113_barrel_shifter_line57;
    wire tmp114_barrel_shifter_line59;
    wire tmp115_barrel_shifter_line59;
    wire[15:0] tmp116_barrel_shifter_line59;
    wire[14:0] tmp117_barrel_shifter_line59;
    wire[15:0] tmp118_barrel_shifter_line59;
    wire[15:0] tmp119_barrel_shifter_line59;
    wire tmp120_barrel_shifter_line62;
    wire tmp121_barrel_shifter_line62;
    wire[31:0] tmp122_barrel_shifter_line62;
    wire[63:0] tmp123_barrel_shifter_line62;
    wire[63:0] tmp124_barrel_shifter_line62;
    wire tmp125_barrel_shifter_line64;
    wire tmp126_barrel_shifter_line64;
    wire[31:0] tmp127_barrel_shifter_line64;
    wire[30:0] tmp128_barrel_shifter_line64;
    wire[31:0] tmp129_barrel_shifter_line64;
    wire[31:0] tmp130_barrel_shifter_line64;
    wire tmp131_barrel_shifter_line69;
    wire tmp132_barrel_shifter_line69;
    wire tmp133_barrel_shifter_line69;
    wire tmp134_barrel_shifter_line69;
    wire tmp135_barrel_shifter_line69;
    wire tmp136_barrel_shifter_line69;
    wire tmp137_barrel_shifter_line69;
    wire tmp138_barrel_shifter_line69;
    wire tmp139_barrel_shifter_line69;
    wire tmp140_barrel_shifter_line69;
    wire tmp141_barrel_shifter_line69;
    wire tmp142_barrel_shifter_line69;
    wire tmp143_barrel_shifter_line69;
    wire tmp144_barrel_shifter_line69;
    wire tmp145_barrel_shifter_line69;
    wire tmp146_barrel_shifter_line69;
    wire tmp147_barrel_shifter_line69;
    wire tmp148_barrel_shifter_line69;
    wire tmp149_barrel_shifter_line69;
    wire tmp150_barrel_shifter_line69;
    wire tmp151_barrel_shifter_line69;
    wire tmp152_barrel_shifter_line69;
    wire tmp153_barrel_shifter_line69;
    wire tmp154_barrel_shifter_line69;
    wire tmp155_barrel_shifter_line69;
    wire tmp156_barrel_shifter_line69;
    wire tmp157_barrel_shifter_line69;
    wire tmp158_barrel_shifter_line69;
    wire tmp159_barrel_shifter_line69;
    wire tmp160_barrel_shifter_line69;
    wire tmp161_barrel_shifter_line69;
    wire tmp162_barrel_shifter_line69;
    wire tmp163_barrel_shifter_line69;
    wire tmp164_barrel_shifter_line69;
    wire tmp165_barrel_shifter_line69;
    wire tmp166_barrel_shifter_line69;
    wire tmp167_barrel_shifter_line69;
    wire tmp168_barrel_shifter_line69;
    wire tmp169_barrel_shifter_line69;
    wire tmp170_barrel_shifter_line69;
    wire tmp171_barrel_shifter_line69;
    wire tmp172_barrel_shifter_line69;
    wire tmp173_barrel_shifter_line69;
    wire tmp174_barrel_shifter_line69;
    wire tmp175_barrel_shifter_line69;
    wire tmp176_barrel_shifter_line69;
    wire tmp177_barrel_shifter_line69;
    wire tmp178_barrel_shifter_line69;
    wire tmp179_barrel_shifter_line69;
    wire tmp180_barrel_shifter_line69;
    wire tmp181_barrel_shifter_line69;
    wire tmp182_barrel_shifter_line69;
    wire tmp183_barrel_shifter_line69;
    wire tmp184_barrel_shifter_line69;
    wire tmp185_barrel_shifter_line69;
    wire tmp186_barrel_shifter_line69;
    wire tmp187_barrel_shifter_line69;
    wire tmp188_barrel_shifter_line69;
    wire tmp189_barrel_shifter_line69;
    wire tmp190_barrel_shifter_line69;
    wire tmp191_barrel_shifter_line69;
    wire tmp192_barrel_shifter_line69;
    wire tmp193_barrel_shifter_line69;
    wire tmp194_barrel_shifter_line69;
    wire tmp195_barrel_shifter_line69;
    wire[63:0] tmp196_barrel_shifter_line69;
    wire[63:0] tmp197_barrel_shifter_line69;
    wire[63:0] tmp198_barrel_shifter_line71;
    wire[63:0] tmp199_barrel_shifter_line71;
    wire[15:0] tmp200_barrel_shifter_line72;
    wire[7:0] tmp201_barrel_shifter_line72;
    wire[3:0] tmp202_barrel_shifter_line72;
    wire[1:0] tmp203_barrel_shifter_line72;
    wire tmp204_barrel_shifter_line72;
    wire tmp205_barrel_shifter_line72;
    wire tmp206_barrel_shifter_line72;
    wire tmp207_barrel_shifter_line72;
    wire tmp208_barrel_shifter_line72;
    wire[1:0] tmp209_barrel_shifter_line72;
    wire tmp210_barrel_shifter_line72;
    wire tmp211_barrel_shifter_line72;
    wire tmp212_barrel_shifter_line72;
    wire tmp213_barrel_shifter_line72;
    wire tmp214_barrel_shifter_line72;
    wire tmp215_barrel_shifter_line72;
    wire[3:0] tmp216_barrel_shifter_line72;
    wire[1:0] tmp217_barrel_shifter_line72;
    wire tmp218_barrel_shifter_line72;
    wire tmp219_barrel_shifter_line72;
    wire tmp220_barrel_shifter_line72;
    wire tmp221_barrel_shifter_line72;
    wire tmp222_barrel_shifter_line72;
    wire[1:0] tmp223_barrel_shifter_line72;
    wire tmp224_barrel_shifter_line72;
    wire tmp225_barrel_shifter_line72;
    wire tmp226_barrel_shifter_line72;
    wire tmp227_barrel_shifter_line72;
    wire tmp228_barrel_shifter_line72;
    wire tmp229_barrel_shifter_line72;
    wire tmp230_barrel_shifter_line72;
    wire[7:0] tmp231_barrel_shifter_line72;
    wire[3:0] tmp232_barrel_shifter_line72;
    wire[1:0] tmp233_barrel_shifter_line72;
    wire tmp234_barrel_shifter_line72;
    wire tmp235_barrel_shifter_line72;
    wire tmp236_barrel_shifter_line72;
    wire tmp237_barrel_shifter_line72;
    wire tmp238_barrel_shifter_line72;
    wire[1:0] tmp239_barrel_shifter_line72;
    wire tmp240_barrel_shifter_line72;
    wire tmp241_barrel_shifter_line72;
    wire tmp242_barrel_shifter_line72;
    wire tmp243_barrel_shifter_line72;
    wire tmp244_barrel_shifter_line72;
    wire tmp245_barrel_shifter_line72;
    wire[3:0] tmp246_barrel_shifter_line72;
    wire[1:0] tmp247_barrel_shifter_line72;
    wire tmp248_barrel_shifter_line72;
    wire tmp249_barrel_shifter_line72;
    wire tmp250_barrel_shifter_line72;
    wire tmp251_barrel_shifter_line72;
    wire tmp252_barrel_shifter_line72;
    wire[1:0] tmp253_barrel_shifter_line72;
    wire tmp254_barrel_shifter_line72;
    wire tmp255_barrel_shifter_line72;
    wire tmp256_barrel_shifter_line72;
    wire tmp257_barrel_shifter_line72;
    wire tmp258_barrel_shifter_line72;
    wire tmp259_barrel_shifter_line72;
    wire tmp260_barrel_shifter_line72;
    wire tmp261_barrel_shifter_line72;
    wire[15:0] tmp262_barrel_shifter_line72;
    wire[7:0] tmp263_barrel_shifter_line72;
    wire[3:0] tmp264_barrel_shifter_line72;
    wire[1:0] tmp265_barrel_shifter_line72;
    wire tmp266_barrel_shifter_line72;
    wire tmp267_barrel_shifter_line72;
    wire tmp268_barrel_shifter_line72;
    wire tmp269_barrel_shifter_line72;
    wire tmp270_barrel_shifter_line72;
    wire[1:0] tmp271_barrel_shifter_line72;
    wire tmp272_barrel_shifter_line72;
    wire tmp273_barrel_shifter_line72;
    wire tmp274_barrel_shifter_line72;
    wire tmp275_barrel_shifter_line72;
    wire tmp276_barrel_shifter_line72;
    wire tmp277_barrel_shifter_line72;
    wire[3:0] tmp278_barrel_shifter_line72;
    wire[1:0] tmp279_barrel_shifter_line72;
    wire tmp280_barrel_shifter_line72;
    wire tmp281_barrel_shifter_line72;
    wire tmp282_barrel_shifter_line72;
    wire tmp283_barrel_shifter_line72;
    wire tmp284_barrel_shifter_line72;
    wire[1:0] tmp285_barrel_shifter_line72;
    wire tmp286_barrel_shifter_line72;
    wire tmp287_barrel_shifter_line72;
    wire tmp288_barrel_shifter_line72;
    wire tmp289_barrel_shifter_line72;
    wire tmp290_barrel_shifter_line72;
    wire tmp291_barrel_shifter_line72;
    wire tmp292_barrel_shifter_line72;
    wire[7:0] tmp293_barrel_shifter_line72;
    wire[3:0] tmp294_barrel_shifter_line72;
    wire[1:0] tmp295_barrel_shifter_line72;
    wire tmp296_barrel_shifter_line72;
    wire tmp297_barrel_shifter_line72;
    wire tmp298_barrel_shifter_line72;
    wire tmp299_barrel_shifter_line72;
    wire tmp300_barrel_shifter_line72;
    wire[1:0] tmp301_barrel_shifter_line72;
    wire tmp302_barrel_shifter_line72;
    wire tmp303_barrel_shifter_line72;
    wire tmp304_barrel_shifter_line72;
    wire tmp305_barrel_shifter_line72;
    wire tmp306_barrel_shifter_line72;
    wire tmp307_barrel_shifter_line72;
    wire[3:0] tmp308_barrel_shifter_line72;
    wire[1:0] tmp309_barrel_shifter_line72;
    wire tmp310_barrel_shifter_line72;
    wire tmp311_barrel_shifter_line72;
    wire tmp312_barrel_shifter_line72;
    wire tmp313_barrel_shifter_line72;
    wire tmp314_barrel_shifter_line72;
    wire[1:0] tmp315_barrel_shifter_line72;
    wire tmp316_barrel_shifter_line72;
    wire tmp317_barrel_shifter_line72;
    wire tmp318_barrel_shifter_line72;
    wire tmp319_barrel_shifter_line72;
    wire tmp320_barrel_shifter_line72;
    wire tmp321_barrel_shifter_line72;
    wire tmp322_barrel_shifter_line72;
    wire tmp323_barrel_shifter_line72;
    wire tmp324_barrel_shifter_line72;
    wire[7:0] tmp325_barrel_shifter_line72;
    wire[3:0] tmp326_barrel_shifter_line72;
    wire[1:0] tmp327_barrel_shifter_line72;
    wire tmp328_barrel_shifter_line72;
    wire tmp329_barrel_shifter_line72;
    wire tmp330_barrel_shifter_line72;
    wire tmp331_barrel_shifter_line72;
    wire tmp332_barrel_shifter_line72;
    wire[1:0] tmp333_barrel_shifter_line72;
    wire tmp334_barrel_shifter_line72;
    wire tmp335_barrel_shifter_line72;
    wire tmp336_barrel_shifter_line72;
    wire tmp337_barrel_shifter_line72;
    wire tmp338_barrel_shifter_line72;
    wire tmp339_barrel_shifter_line72;
    wire[3:0] tmp340_barrel_shifter_line72;
    wire[1:0] tmp341_barrel_shifter_line72;
    wire tmp342_barrel_shifter_line72;
    wire tmp343_barrel_shifter_line72;
    wire tmp344_barrel_shifter_line72;
    wire tmp345_barrel_shifter_line72;
    wire tmp346_barrel_shifter_line72;
    wire[1:0] tmp347_barrel_shifter_line72;
    wire tmp348_barrel_shifter_line72;
    wire tmp349_barrel_shifter_line72;
    wire tmp350_barrel_shifter_line72;
    wire tmp351_barrel_shifter_line72;
    wire tmp352_barrel_shifter_line72;
    wire tmp353_barrel_shifter_line72;
    wire tmp354_barrel_shifter_line72;
    wire[7:0] tmp355_barrel_shifter_line72;
    wire[3:0] tmp356_barrel_shifter_line72;
    wire[1:0] tmp357_barrel_shifter_line72;
    wire tmp358_barrel_shifter_line72;
    wire tmp359_barrel_shifter_line72;
    wire tmp360_barrel_shifter_line72;
    wire tmp361_barrel_shifter_line72;
    wire tmp362_barrel_shifter_line72;
    wire[1:0] tmp363_barrel_shifter_line72;
    wire tmp364_barrel_shifter_line72;
    wire tmp365_barrel_shifter_line72;
    wire tmp366_barrel_shifter_line72;
    wire tmp367_barrel_shifter_line72;
    wire tmp368_barrel_shifter_line72;
    wire tmp369_barrel_shifter_line72;
    wire[3:0] tmp370_barrel_shifter_line72;
    wire[1:0] tmp371_barrel_shifter_line72;
    wire tmp372_barrel_shifter_line72;
    wire tmp373_barrel_shifter_line72;
    wire tmp374_barrel_shifter_line72;
    wire tmp375_barrel_shifter_line72;
    wire tmp376_barrel_shifter_line72;
    wire[1:0] tmp377_barrel_shifter_line72;
    wire tmp378_barrel_shifter_line72;
    wire tmp379_barrel_shifter_line72;
    wire tmp380_barrel_shifter_line72;
    wire tmp381_barrel_shifter_line72;
    wire tmp382_barrel_shifter_line72;
    wire tmp383_barrel_shifter_line72;
    wire tmp384_barrel_shifter_line72;
    wire tmp385_barrel_shifter_line72;
    wire tmp386_barrel_shifter_line72;
    wire[3:0] tmp387_barrel_shifter_line72;
    wire[1:0] tmp388_barrel_shifter_line72;
    wire tmp389_barrel_shifter_line72;
    wire tmp390_barrel_shifter_line72;
    wire tmp391_barrel_shifter_line72;
    wire tmp392_barrel_shifter_line72;
    wire tmp393_barrel_shifter_line72;
    wire[1:0] tmp394_barrel_shifter_line72;
    wire tmp395_barrel_shifter_line72;
    wire tmp396_barrel_shifter_line72;
    wire tmp397_barrel_shifter_line72;
    wire tmp398_barrel_shifter_line72;
    wire tmp399_barrel_shifter_line72;
    wire tmp400_barrel_shifter_line72;
    wire[3:0] tmp401_barrel_shifter_line72;
    wire[1:0] tmp402_barrel_shifter_line72;
    wire tmp403_barrel_shifter_line72;
    wire tmp404_barrel_shifter_line72;
    wire tmp405_barrel_shifter_line72;
    wire tmp406_barrel_shifter_line72;
    wire tmp407_barrel_shifter_line72;
    wire[1:0] tmp408_barrel_shifter_line72;
    wire tmp409_barrel_shifter_line72;
    wire tmp410_barrel_shifter_line72;
    wire tmp411_barrel_shifter_line72;
    wire tmp412_barrel_shifter_line72;
    wire tmp413_barrel_shifter_line72;
    wire tmp414_barrel_shifter_line72;
    wire tmp415_barrel_shifter_line72;
    wire tmp416_barrel_shifter_line72;
    wire[1:0] tmp417_barrel_shifter_line72;
    wire tmp418_barrel_shifter_line72;
    wire tmp419_barrel_shifter_line72;
    wire tmp420_barrel_shifter_line72;
    wire tmp421_barrel_shifter_line72;
    wire tmp422_barrel_shifter_line72;
    wire[1:0] tmp423_barrel_shifter_line72;
    wire tmp424_barrel_shifter_line72;
    wire tmp425_barrel_shifter_line72;
    wire tmp426_barrel_shifter_line72;
    wire tmp427_barrel_shifter_line72;
    wire tmp428_barrel_shifter_line72;
    wire tmp429_barrel_shifter_line72;
    wire tmp430_barrel_shifter_line72;
    wire tmp431_barrel_shifter_line72;
    wire tmp432_barrel_shifter_line72;
    wire tmp433_barrel_shifter_line72;
    wire tmp434_barrel_shifter_line72;
    wire tmp435_barrel_shifter_line72;
    wire tmp436_barrel_shifter_line72;
    wire tmp437_barrel_shifter_line72;
    wire tmp438_barrel_shifter_line72;

    // Combinational
    assign const_0_0 = 0;
    assign const_1_0 = 0;
    assign const_2_0 = 0;
    assign const_3_0 = 0;
    assign const_4_0 = 0;
    assign const_5_0 = 0;
    assign const_6_0 = 0;
    assign const_7_0 = 0;
    assign const_8_0 = 0;
    assign const_9_0 = 0;
    assign const_10_0 = 0;
    assign const_11_0 = 0;
    assign const_12_0 = 0;
    assign const_13_0 = 0;
    assign const_14_0 = 0;
    assign const_15_0 = 0;
    assign const_16_0 = 0;
    assign const_17_0 = 0;
    assign const_18_0 = 0;
    assign const_19_0 = 0;
    assign const_20_0 = 0;
    assign const_21_0 = 0;
    assign const_22_0 = 0;
    assign const_23_0 = 0;
    assign const_24_0 = 0;
    assign overflow = tmp438_barrel_shifter_line72;
    assign reverse_in = tmp66_barrel_shifter_line25;
    assign reverse_out = tmp197_barrel_shifter_line69;
    assign s = tmp199_barrel_shifter_line71;
    assign shift_1 = tmp71_barrel_shifter_line37;
    assign shift_2 = tmp80_barrel_shifter_line42;
    assign shift_4 = tmp91_barrel_shifter_line47;
    assign shift_8 = tmp102_barrel_shifter_line52;
    assign shift_16 = tmp113_barrel_shifter_line57;
    assign shift_32 = tmp124_barrel_shifter_line62;
    assign shift_off_1 = tmp75_barrel_shifter_line39;
    assign shift_off_2 = tmp86_barrel_shifter_line44;
    assign shift_off_4 = tmp97_barrel_shifter_line49;
    assign shift_off_8 = tmp108_barrel_shifter_line54;
    assign shift_off_16 = tmp119_barrel_shifter_line59;
    assign shift_off_32 = tmp130_barrel_shifter_line64;
    assign tmp0_barrel_shifter_line25 = direction == const_0_0;
    assign tmp1_barrel_shifter_line25 = {a[63]};
    assign tmp2_barrel_shifter_line25 = {a[62]};
    assign tmp3_barrel_shifter_line25 = {a[61]};
    assign tmp4_barrel_shifter_line25 = {a[60]};
    assign tmp5_barrel_shifter_line25 = {a[59]};
    assign tmp6_barrel_shifter_line25 = {a[58]};
    assign tmp7_barrel_shifter_line25 = {a[57]};
    assign tmp8_barrel_shifter_line25 = {a[56]};
    assign tmp9_barrel_shifter_line25 = {a[55]};
    assign tmp10_barrel_shifter_line25 = {a[54]};
    assign tmp11_barrel_shifter_line25 = {a[53]};
    assign tmp12_barrel_shifter_line25 = {a[52]};
    assign tmp13_barrel_shifter_line25 = {a[51]};
    assign tmp14_barrel_shifter_line25 = {a[50]};
    assign tmp15_barrel_shifter_line25 = {a[49]};
    assign tmp16_barrel_shifter_line25 = {a[48]};
    assign tmp17_barrel_shifter_line25 = {a[47]};
    assign tmp18_barrel_shifter_line25 = {a[46]};
    assign tmp19_barrel_shifter_line25 = {a[45]};
    assign tmp20_barrel_shifter_line25 = {a[44]};
    assign tmp21_barrel_shifter_line25 = {a[43]};
    assign tmp22_barrel_shifter_line25 = {a[42]};
    assign tmp23_barrel_shifter_line25 = {a[41]};
    assign tmp24_barrel_shifter_line25 = {a[40]};
    assign tmp25_barrel_shifter_line25 = {a[39]};
    assign tmp26_barrel_shifter_line25 = {a[38]};
    assign tmp27_barrel_shifter_line25 = {a[37]};
    assign tmp28_barrel_shifter_line25 = {a[36]};
    assign tmp29_barrel_shifter_line25 = {a[35]};
    assign tmp30_barrel_shifter_line25 = {a[34]};
    assign tmp31_barrel_shifter_line25 = {a[33]};
    assign tmp32_barrel_shifter_line25 = {a[32]};
    assign tmp33_barrel_shifter_line25 = {a[31]};
    assign tmp34_barrel_shifter_line25 = {a[30]};
    assign tmp35_barrel_shifter_line25 = {a[29]};
    assign tmp36_barrel_shifter_line25 = {a[28]};
    assign tmp37_barrel_shifter_line25 = {a[27]};
    assign tmp38_barrel_shifter_line25 = {a[26]};
    assign tmp39_barrel_shifter_line25 = {a[25]};
    assign tmp40_barrel_shifter_line25 = {a[24]};
    assign tmp41_barrel_shifter_line25 = {a[23]};
    assign tmp42_barrel_shifter_line25 = {a[22]};
    assign tmp43_barrel_shifter_line25 = {a[21]};
    assign tmp44_barrel_shifter_line25 = {a[20]};
    assign tmp45_barrel_shifter_line25 = {a[19]};
    assign tmp46_barrel_shifter_line25 = {a[18]};
    assign tmp47_barrel_shifter_line25 = {a[17]};
    assign tmp48_barrel_shifter_line25 = {a[16]};
    assign tmp49_barrel_shifter_line25 = {a[15]};
    assign tmp50_barrel_shifter_line25 = {a[14]};
    assign tmp51_barrel_shifter_line25 = {a[13]};
    assign tmp52_barrel_shifter_line25 = {a[12]};
    assign tmp53_barrel_shifter_line25 = {a[11]};
    assign tmp54_barrel_shifter_line25 = {a[10]};
    assign tmp55_barrel_shifter_line25 = {a[9]};
    assign tmp56_barrel_shifter_line25 = {a[8]};
    assign tmp57_barrel_shifter_line25 = {a[7]};
    assign tmp58_barrel_shifter_line25 = {a[6]};
    assign tmp59_barrel_shifter_line25 = {a[5]};
    assign tmp60_barrel_shifter_line25 = {a[4]};
    assign tmp61_barrel_shifter_line25 = {a[3]};
    assign tmp62_barrel_shifter_line25 = {a[2]};
    assign tmp63_barrel_shifter_line25 = {a[1]};
    assign tmp64_barrel_shifter_line25 = {a[0]};
    assign tmp65_barrel_shifter_line25 = {tmp64_barrel_shifter_line25, tmp63_barrel_shifter_line25, tmp62_barrel_shifter_line25, tmp61_barrel_shifter_line25, tmp60_barrel_shifter_line25, tmp59_barrel_shifter_line25, tmp58_barrel_shifter_line25, tmp57_barrel_shifter_line25, tmp56_barrel_shifter_line25, tmp55_barrel_shifter_line25, tmp54_barrel_shifter_line25, tmp53_barrel_shifter_line25, tmp52_barrel_shifter_line25, tmp51_barrel_shifter_line25, tmp50_barrel_shifter_line25, tmp49_barrel_shifter_line25, tmp48_barrel_shifter_line25, tmp47_barrel_shifter_line25, tmp46_barrel_shifter_line25, tmp45_barrel_shifter_line25, tmp44_barrel_shifter_line25, tmp43_barrel_shifter_line25, tmp42_barrel_shifter_line25, tmp41_barrel_shifter_line25, tmp40_barrel_shifter_line25, tmp39_barrel_shifter_line25, tmp38_barrel_shifter_line25, tmp37_barrel_shifter_line25, tmp36_barrel_shifter_line25, tmp35_barrel_shifter_line25, tmp34_barrel_shifter_line25, tmp33_barrel_shifter_line25, tmp32_barrel_shifter_line25, tmp31_barrel_shifter_line25, tmp30_barrel_shifter_line25, tmp29_barrel_shifter_line25, tmp28_barrel_shifter_line25, tmp27_barrel_shifter_line25, tmp26_barrel_shifter_line25, tmp25_barrel_shifter_line25, tmp24_barrel_shifter_line25, tmp23_barrel_shifter_line25, tmp22_barrel_shifter_line25, tmp21_barrel_shifter_line25, tmp20_barrel_shifter_line25, tmp19_barrel_shifter_line25, tmp18_barrel_shifter_line25, tmp17_barrel_shifter_line25, tmp16_barrel_shifter_line25, tmp15_barrel_shifter_line25, tmp14_barrel_shifter_line25, tmp13_barrel_shifter_line25, tmp12_barrel_shifter_line25, tmp11_barrel_shifter_line25, tmp10_barrel_shifter_line25, tmp9_barrel_shifter_line25, tmp8_barrel_shifter_line25, tmp7_barrel_shifter_line25, tmp6_barrel_shifter_line25, tmp5_barrel_shifter_line25, tmp4_barrel_shifter_line25, tmp3_barrel_shifter_line25, tmp2_barrel_shifter_line25, tmp1_barrel_shifter_line25};
    assign tmp66_barrel_shifter_line25 = tmp0_barrel_shifter_line25 ? a : tmp65_barrel_shifter_line25;
    assign tmp67_barrel_shifter_line37 = {n[0]};
    assign tmp68_barrel_shifter_line37 = tmp67_barrel_shifter_line37 == const_1_0;
    assign tmp69_barrel_shifter_line37 = {reverse_in[62], reverse_in[61], reverse_in[60], reverse_in[59], reverse_in[58], reverse_in[57], reverse_in[56], reverse_in[55], reverse_in[54], reverse_in[53], reverse_in[52], reverse_in[51], reverse_in[50], reverse_in[49], reverse_in[48], reverse_in[47], reverse_in[46], reverse_in[45], reverse_in[44], reverse_in[43], reverse_in[42], reverse_in[41], reverse_in[40], reverse_in[39], reverse_in[38], reverse_in[37], reverse_in[36], reverse_in[35], reverse_in[34], reverse_in[33], reverse_in[32], reverse_in[31], reverse_in[30], reverse_in[29], reverse_in[28], reverse_in[27], reverse_in[26], reverse_in[25], reverse_in[24], reverse_in[23], reverse_in[22], reverse_in[21], reverse_in[20], reverse_in[19], reverse_in[18], reverse_in[17], reverse_in[16], reverse_in[15], reverse_in[14], reverse_in[13], reverse_in[12], reverse_in[11], reverse_in[10], reverse_in[9], reverse_in[8], reverse_in[7], reverse_in[6], reverse_in[5], reverse_in[4], reverse_in[3], reverse_in[2], reverse_in[1], reverse_in[0]};
    assign tmp70_barrel_shifter_line37 = {tmp69_barrel_shifter_line37, shift_in};
    assign tmp71_barrel_shifter_line37 = tmp68_barrel_shifter_line37 ? reverse_in : tmp70_barrel_shifter_line37;
    assign tmp72_barrel_shifter_line39 = {n[0]};
    assign tmp73_barrel_shifter_line39 = tmp72_barrel_shifter_line39 == const_2_0;
    assign tmp74_barrel_shifter_line39 = {reverse_in[63]};
    assign tmp75_barrel_shifter_line39 = tmp73_barrel_shifter_line39 ? const_3_0 : tmp74_barrel_shifter_line39;
    assign tmp76_barrel_shifter_line42 = {n[1]};
    assign tmp77_barrel_shifter_line42 = tmp76_barrel_shifter_line42 == const_4_0;
    assign tmp78_barrel_shifter_line42 = {shift_1[61], shift_1[60], shift_1[59], shift_1[58], shift_1[57], shift_1[56], shift_1[55], shift_1[54], shift_1[53], shift_1[52], shift_1[51], shift_1[50], shift_1[49], shift_1[48], shift_1[47], shift_1[46], shift_1[45], shift_1[44], shift_1[43], shift_1[42], shift_1[41], shift_1[40], shift_1[39], shift_1[38], shift_1[37], shift_1[36], shift_1[35], shift_1[34], shift_1[33], shift_1[32], shift_1[31], shift_1[30], shift_1[29], shift_1[28], shift_1[27], shift_1[26], shift_1[25], shift_1[24], shift_1[23], shift_1[22], shift_1[21], shift_1[20], shift_1[19], shift_1[18], shift_1[17], shift_1[16], shift_1[15], shift_1[14], shift_1[13], shift_1[12], shift_1[11], shift_1[10], shift_1[9], shift_1[8], shift_1[7], shift_1[6], shift_1[5], shift_1[4], shift_1[3], shift_1[2], shift_1[1], shift_1[0]};
    assign tmp79_barrel_shifter_line42 = {tmp78_barrel_shifter_line42, shift_in, shift_in};
    assign tmp80_barrel_shifter_line42 = tmp77_barrel_shifter_line42 ? shift_1 : tmp79_barrel_shifter_line42;
    assign tmp81_barrel_shifter_line44 = {n[1]};
    assign tmp82_barrel_shifter_line44 = tmp81_barrel_shifter_line44 == const_5_0;
    assign tmp83_barrel_shifter_line44 = {shift_1[63], shift_1[62]};
    assign tmp84_barrel_shifter_line44 = {const_7_0};
    assign tmp85_barrel_shifter_line44 = {tmp84_barrel_shifter_line44, const_6_0};
    assign tmp86_barrel_shifter_line44 = tmp82_barrel_shifter_line44 ? tmp85_barrel_shifter_line44 : tmp83_barrel_shifter_line44;
    assign tmp87_barrel_shifter_line47 = {n[2]};
    assign tmp88_barrel_shifter_line47 = tmp87_barrel_shifter_line47 == const_8_0;
    assign tmp89_barrel_shifter_line47 = {shift_2[59], shift_2[58], shift_2[57], shift_2[56], shift_2[55], shift_2[54], shift_2[53], shift_2[52], shift_2[51], shift_2[50], shift_2[49], shift_2[48], shift_2[47], shift_2[46], shift_2[45], shift_2[44], shift_2[43], shift_2[42], shift_2[41], shift_2[40], shift_2[39], shift_2[38], shift_2[37], shift_2[36], shift_2[35], shift_2[34], shift_2[33], shift_2[32], shift_2[31], shift_2[30], shift_2[29], shift_2[28], shift_2[27], shift_2[26], shift_2[25], shift_2[24], shift_2[23], shift_2[22], shift_2[21], shift_2[20], shift_2[19], shift_2[18], shift_2[17], shift_2[16], shift_2[15], shift_2[14], shift_2[13], shift_2[12], shift_2[11], shift_2[10], shift_2[9], shift_2[8], shift_2[7], shift_2[6], shift_2[5], shift_2[4], shift_2[3], shift_2[2], shift_2[1], shift_2[0]};
    assign tmp90_barrel_shifter_line47 = {tmp89_barrel_shifter_line47, shift_in, shift_in, shift_in, shift_in};
    assign tmp91_barrel_shifter_line47 = tmp88_barrel_shifter_line47 ? shift_2 : tmp90_barrel_shifter_line47;
    assign tmp92_barrel_shifter_line49 = {n[1]};
    assign tmp93_barrel_shifter_line49 = tmp92_barrel_shifter_line49 == const_9_0;
    assign tmp94_barrel_shifter_line49 = {shift_2[63], shift_2[62], shift_2[61], shift_2[60]};
    assign tmp95_barrel_shifter_line49 = {const_11_0, const_11_0, const_11_0};
    assign tmp96_barrel_shifter_line49 = {tmp95_barrel_shifter_line49, const_10_0};
    assign tmp97_barrel_shifter_line49 = tmp93_barrel_shifter_line49 ? tmp96_barrel_shifter_line49 : tmp94_barrel_shifter_line49;
    assign tmp98_barrel_shifter_line52 = {n[3]};
    assign tmp99_barrel_shifter_line52 = tmp98_barrel_shifter_line52 == const_12_0;
    assign tmp100_barrel_shifter_line52 = {shift_4[55], shift_4[54], shift_4[53], shift_4[52], shift_4[51], shift_4[50], shift_4[49], shift_4[48], shift_4[47], shift_4[46], shift_4[45], shift_4[44], shift_4[43], shift_4[42], shift_4[41], shift_4[40], shift_4[39], shift_4[38], shift_4[37], shift_4[36], shift_4[35], shift_4[34], shift_4[33], shift_4[32], shift_4[31], shift_4[30], shift_4[29], shift_4[28], shift_4[27], shift_4[26], shift_4[25], shift_4[24], shift_4[23], shift_4[22], shift_4[21], shift_4[20], shift_4[19], shift_4[18], shift_4[17], shift_4[16], shift_4[15], shift_4[14], shift_4[13], shift_4[12], shift_4[11], shift_4[10], shift_4[9], shift_4[8], shift_4[7], shift_4[6], shift_4[5], shift_4[4], shift_4[3], shift_4[2], shift_4[1], shift_4[0]};
    assign tmp101_barrel_shifter_line52 = {tmp100_barrel_shifter_line52, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in};
    assign tmp102_barrel_shifter_line52 = tmp99_barrel_shifter_line52 ? shift_4 : tmp101_barrel_shifter_line52;
    assign tmp103_barrel_shifter_line54 = {n[1]};
    assign tmp104_barrel_shifter_line54 = tmp103_barrel_shifter_line54 == const_13_0;
    assign tmp105_barrel_shifter_line54 = {shift_4[63], shift_4[62], shift_4[61], shift_4[60], shift_4[59], shift_4[58], shift_4[57], shift_4[56]};
    assign tmp106_barrel_shifter_line54 = {const_15_0, const_15_0, const_15_0, const_15_0, const_15_0, const_15_0, const_15_0};
    assign tmp107_barrel_shifter_line54 = {tmp106_barrel_shifter_line54, const_14_0};
    assign tmp108_barrel_shifter_line54 = tmp104_barrel_shifter_line54 ? tmp107_barrel_shifter_line54 : tmp105_barrel_shifter_line54;
    assign tmp109_barrel_shifter_line57 = {n[4]};
    assign tmp110_barrel_shifter_line57 = tmp109_barrel_shifter_line57 == const_16_0;
    assign tmp111_barrel_shifter_line57 = {shift_8[47], shift_8[46], shift_8[45], shift_8[44], shift_8[43], shift_8[42], shift_8[41], shift_8[40], shift_8[39], shift_8[38], shift_8[37], shift_8[36], shift_8[35], shift_8[34], shift_8[33], shift_8[32], shift_8[31], shift_8[30], shift_8[29], shift_8[28], shift_8[27], shift_8[26], shift_8[25], shift_8[24], shift_8[23], shift_8[22], shift_8[21], shift_8[20], shift_8[19], shift_8[18], shift_8[17], shift_8[16], shift_8[15], shift_8[14], shift_8[13], shift_8[12], shift_8[11], shift_8[10], shift_8[9], shift_8[8], shift_8[7], shift_8[6], shift_8[5], shift_8[4], shift_8[3], shift_8[2], shift_8[1], shift_8[0]};
    assign tmp112_barrel_shifter_line57 = {tmp111_barrel_shifter_line57, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in};
    assign tmp113_barrel_shifter_line57 = tmp110_barrel_shifter_line57 ? shift_8 : tmp112_barrel_shifter_line57;
    assign tmp114_barrel_shifter_line59 = {n[1]};
    assign tmp115_barrel_shifter_line59 = tmp114_barrel_shifter_line59 == const_17_0;
    assign tmp116_barrel_shifter_line59 = {shift_8[63], shift_8[62], shift_8[61], shift_8[60], shift_8[59], shift_8[58], shift_8[57], shift_8[56], shift_8[55], shift_8[54], shift_8[53], shift_8[52], shift_8[51], shift_8[50], shift_8[49], shift_8[48]};
    assign tmp117_barrel_shifter_line59 = {const_19_0, const_19_0, const_19_0, const_19_0, const_19_0, const_19_0, const_19_0, const_19_0, const_19_0, const_19_0, const_19_0, const_19_0, const_19_0, const_19_0, const_19_0};
    assign tmp118_barrel_shifter_line59 = {tmp117_barrel_shifter_line59, const_18_0};
    assign tmp119_barrel_shifter_line59 = tmp115_barrel_shifter_line59 ? tmp118_barrel_shifter_line59 : tmp116_barrel_shifter_line59;
    assign tmp120_barrel_shifter_line62 = {n[5]};
    assign tmp121_barrel_shifter_line62 = tmp120_barrel_shifter_line62 == const_20_0;
    assign tmp122_barrel_shifter_line62 = {shift_16[31], shift_16[30], shift_16[29], shift_16[28], shift_16[27], shift_16[26], shift_16[25], shift_16[24], shift_16[23], shift_16[22], shift_16[21], shift_16[20], shift_16[19], shift_16[18], shift_16[17], shift_16[16], shift_16[15], shift_16[14], shift_16[13], shift_16[12], shift_16[11], shift_16[10], shift_16[9], shift_16[8], shift_16[7], shift_16[6], shift_16[5], shift_16[4], shift_16[3], shift_16[2], shift_16[1], shift_16[0]};
    assign tmp123_barrel_shifter_line62 = {tmp122_barrel_shifter_line62, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in};
    assign tmp124_barrel_shifter_line62 = tmp121_barrel_shifter_line62 ? shift_16 : tmp123_barrel_shifter_line62;
    assign tmp125_barrel_shifter_line64 = {n[1]};
    assign tmp126_barrel_shifter_line64 = tmp125_barrel_shifter_line64 == const_21_0;
    assign tmp127_barrel_shifter_line64 = {shift_16[63], shift_16[62], shift_16[61], shift_16[60], shift_16[59], shift_16[58], shift_16[57], shift_16[56], shift_16[55], shift_16[54], shift_16[53], shift_16[52], shift_16[51], shift_16[50], shift_16[49], shift_16[48], shift_16[47], shift_16[46], shift_16[45], shift_16[44], shift_16[43], shift_16[42], shift_16[41], shift_16[40], shift_16[39], shift_16[38], shift_16[37], shift_16[36], shift_16[35], shift_16[34], shift_16[33], shift_16[32]};
    assign tmp128_barrel_shifter_line64 = {const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0, const_23_0};
    assign tmp129_barrel_shifter_line64 = {tmp128_barrel_shifter_line64, const_22_0};
    assign tmp130_barrel_shifter_line64 = tmp126_barrel_shifter_line64 ? tmp129_barrel_shifter_line64 : tmp127_barrel_shifter_line64;
    assign tmp131_barrel_shifter_line69 = direction == const_24_0;
    assign tmp132_barrel_shifter_line69 = {shift_32[63]};
    assign tmp133_barrel_shifter_line69 = {shift_32[62]};
    assign tmp134_barrel_shifter_line69 = {shift_32[61]};
    assign tmp135_barrel_shifter_line69 = {shift_32[60]};
    assign tmp136_barrel_shifter_line69 = {shift_32[59]};
    assign tmp137_barrel_shifter_line69 = {shift_32[58]};
    assign tmp138_barrel_shifter_line69 = {shift_32[57]};
    assign tmp139_barrel_shifter_line69 = {shift_32[56]};
    assign tmp140_barrel_shifter_line69 = {shift_32[55]};
    assign tmp141_barrel_shifter_line69 = {shift_32[54]};
    assign tmp142_barrel_shifter_line69 = {shift_32[53]};
    assign tmp143_barrel_shifter_line69 = {shift_32[52]};
    assign tmp144_barrel_shifter_line69 = {shift_32[51]};
    assign tmp145_barrel_shifter_line69 = {shift_32[50]};
    assign tmp146_barrel_shifter_line69 = {shift_32[49]};
    assign tmp147_barrel_shifter_line69 = {shift_32[48]};
    assign tmp148_barrel_shifter_line69 = {shift_32[47]};
    assign tmp149_barrel_shifter_line69 = {shift_32[46]};
    assign tmp150_barrel_shifter_line69 = {shift_32[45]};
    assign tmp151_barrel_shifter_line69 = {shift_32[44]};
    assign tmp152_barrel_shifter_line69 = {shift_32[43]};
    assign tmp153_barrel_shifter_line69 = {shift_32[42]};
    assign tmp154_barrel_shifter_line69 = {shift_32[41]};
    assign tmp155_barrel_shifter_line69 = {shift_32[40]};
    assign tmp156_barrel_shifter_line69 = {shift_32[39]};
    assign tmp157_barrel_shifter_line69 = {shift_32[38]};
    assign tmp158_barrel_shifter_line69 = {shift_32[37]};
    assign tmp159_barrel_shifter_line69 = {shift_32[36]};
    assign tmp160_barrel_shifter_line69 = {shift_32[35]};
    assign tmp161_barrel_shifter_line69 = {shift_32[34]};
    assign tmp162_barrel_shifter_line69 = {shift_32[33]};
    assign tmp163_barrel_shifter_line69 = {shift_32[32]};
    assign tmp164_barrel_shifter_line69 = {shift_32[31]};
    assign tmp165_barrel_shifter_line69 = {shift_32[30]};
    assign tmp166_barrel_shifter_line69 = {shift_32[29]};
    assign tmp167_barrel_shifter_line69 = {shift_32[28]};
    assign tmp168_barrel_shifter_line69 = {shift_32[27]};
    assign tmp169_barrel_shifter_line69 = {shift_32[26]};
    assign tmp170_barrel_shifter_line69 = {shift_32[25]};
    assign tmp171_barrel_shifter_line69 = {shift_32[24]};
    assign tmp172_barrel_shifter_line69 = {shift_32[23]};
    assign tmp173_barrel_shifter_line69 = {shift_32[22]};
    assign tmp174_barrel_shifter_line69 = {shift_32[21]};
    assign tmp175_barrel_shifter_line69 = {shift_32[20]};
    assign tmp176_barrel_shifter_line69 = {shift_32[19]};
    assign tmp177_barrel_shifter_line69 = {shift_32[18]};
    assign tmp178_barrel_shifter_line69 = {shift_32[17]};
    assign tmp179_barrel_shifter_line69 = {shift_32[16]};
    assign tmp180_barrel_shifter_line69 = {shift_32[15]};
    assign tmp181_barrel_shifter_line69 = {shift_32[14]};
    assign tmp182_barrel_shifter_line69 = {shift_32[13]};
    assign tmp183_barrel_shifter_line69 = {shift_32[12]};
    assign tmp184_barrel_shifter_line69 = {shift_32[11]};
    assign tmp185_barrel_shifter_line69 = {shift_32[10]};
    assign tmp186_barrel_shifter_line69 = {shift_32[9]};
    assign tmp187_barrel_shifter_line69 = {shift_32[8]};
    assign tmp188_barrel_shifter_line69 = {shift_32[7]};
    assign tmp189_barrel_shifter_line69 = {shift_32[6]};
    assign tmp190_barrel_shifter_line69 = {shift_32[5]};
    assign tmp191_barrel_shifter_line69 = {shift_32[4]};
    assign tmp192_barrel_shifter_line69 = {shift_32[3]};
    assign tmp193_barrel_shifter_line69 = {shift_32[2]};
    assign tmp194_barrel_shifter_line69 = {shift_32[1]};
    assign tmp195_barrel_shifter_line69 = {shift_32[0]};
    assign tmp196_barrel_shifter_line69 = {tmp195_barrel_shifter_line69, tmp194_barrel_shifter_line69, tmp193_barrel_shifter_line69, tmp192_barrel_shifter_line69, tmp191_barrel_shifter_line69, tmp190_barrel_shifter_line69, tmp189_barrel_shifter_line69, tmp188_barrel_shifter_line69, tmp187_barrel_shifter_line69, tmp186_barrel_shifter_line69, tmp185_barrel_shifter_line69, tmp184_barrel_shifter_line69, tmp183_barrel_shifter_line69, tmp182_barrel_shifter_line69, tmp181_barrel_shifter_line69, tmp180_barrel_shifter_line69, tmp179_barrel_shifter_line69, tmp178_barrel_shifter_line69, tmp177_barrel_shifter_line69, tmp176_barrel_shifter_line69, tmp175_barrel_shifter_line69, tmp174_barrel_shifter_line69, tmp173_barrel_shifter_line69, tmp172_barrel_shifter_line69, tmp171_barrel_shifter_line69, tmp170_barrel_shifter_line69, tmp169_barrel_shifter_line69, tmp168_barrel_shifter_line69, tmp167_barrel_shifter_line69, tmp166_barrel_shifter_line69, tmp165_barrel_shifter_line69, tmp164_barrel_shifter_line69, tmp163_barrel_shifter_line69, tmp162_barrel_shifter_line69, tmp161_barrel_shifter_line69, tmp160_barrel_shifter_line69, tmp159_barrel_shifter_line69, tmp158_barrel_shifter_line69, tmp157_barrel_shifter_line69, tmp156_barrel_shifter_line69, tmp155_barrel_shifter_line69, tmp154_barrel_shifter_line69, tmp153_barrel_shifter_line69, tmp152_barrel_shifter_line69, tmp151_barrel_shifter_line69, tmp150_barrel_shifter_line69, tmp149_barrel_shifter_line69, tmp148_barrel_shifter_line69, tmp147_barrel_shifter_line69, tmp146_barrel_shifter_line69, tmp145_barrel_shifter_line69, tmp144_barrel_shifter_line69, tmp143_barrel_shifter_line69, tmp142_barrel_shifter_line69, tmp141_barrel_shifter_line69, tmp140_barrel_shifter_line69, tmp139_barrel_shifter_line69, tmp138_barrel_shifter_line69, tmp137_barrel_shifter_line69, tmp136_barrel_shifter_line69, tmp135_barrel_shifter_line69, tmp134_barrel_shifter_line69, tmp133_barrel_shifter_line69, tmp132_barrel_shifter_line69};
    assign tmp197_barrel_shifter_line69 = tmp131_barrel_shifter_line69 ? shift_32 : tmp196_barrel_shifter_line69;
    assign tmp198_barrel_shifter_line71 = ~reverse_out;
    assign tmp199_barrel_shifter_line71 = invert ? tmp198_barrel_shifter_line71 : reverse_out;
    assign tmp200_barrel_shifter_line72 = {shift_off_32[15], shift_off_32[14], shift_off_32[13], shift_off_32[12], shift_off_32[11], shift_off_32[10], shift_off_32[9], shift_off_32[8], shift_off_32[7], shift_off_32[6], shift_off_32[5], shift_off_32[4], shift_off_32[3], shift_off_32[2], shift_off_32[1], shift_off_32[0]};
    assign tmp201_barrel_shifter_line72 = {tmp200_barrel_shifter_line72[7], tmp200_barrel_shifter_line72[6], tmp200_barrel_shifter_line72[5], tmp200_barrel_shifter_line72[4], tmp200_barrel_shifter_line72[3], tmp200_barrel_shifter_line72[2], tmp200_barrel_shifter_line72[1], tmp200_barrel_shifter_line72[0]};
    assign tmp202_barrel_shifter_line72 = {tmp201_barrel_shifter_line72[3], tmp201_barrel_shifter_line72[2], tmp201_barrel_shifter_line72[1], tmp201_barrel_shifter_line72[0]};
    assign tmp203_barrel_shifter_line72 = {tmp202_barrel_shifter_line72[1], tmp202_barrel_shifter_line72[0]};
    assign tmp204_barrel_shifter_line72 = {tmp203_barrel_shifter_line72[0]};
    assign tmp205_barrel_shifter_line72 = {tmp204_barrel_shifter_line72};
    assign tmp206_barrel_shifter_line72 = {tmp203_barrel_shifter_line72[1]};
    assign tmp207_barrel_shifter_line72 = {tmp206_barrel_shifter_line72};
    assign tmp208_barrel_shifter_line72 = tmp205_barrel_shifter_line72 | tmp207_barrel_shifter_line72;
    assign tmp209_barrel_shifter_line72 = {tmp202_barrel_shifter_line72[3], tmp202_barrel_shifter_line72[2]};
    assign tmp210_barrel_shifter_line72 = {tmp209_barrel_shifter_line72[0]};
    assign tmp211_barrel_shifter_line72 = {tmp210_barrel_shifter_line72};
    assign tmp212_barrel_shifter_line72 = {tmp209_barrel_shifter_line72[1]};
    assign tmp213_barrel_shifter_line72 = {tmp212_barrel_shifter_line72};
    assign tmp214_barrel_shifter_line72 = tmp211_barrel_shifter_line72 | tmp213_barrel_shifter_line72;
    assign tmp215_barrel_shifter_line72 = tmp208_barrel_shifter_line72 | tmp214_barrel_shifter_line72;
    assign tmp216_barrel_shifter_line72 = {tmp201_barrel_shifter_line72[7], tmp201_barrel_shifter_line72[6], tmp201_barrel_shifter_line72[5], tmp201_barrel_shifter_line72[4]};
    assign tmp217_barrel_shifter_line72 = {tmp216_barrel_shifter_line72[1], tmp216_barrel_shifter_line72[0]};
    assign tmp218_barrel_shifter_line72 = {tmp217_barrel_shifter_line72[0]};
    assign tmp219_barrel_shifter_line72 = {tmp218_barrel_shifter_line72};
    assign tmp220_barrel_shifter_line72 = {tmp217_barrel_shifter_line72[1]};
    assign tmp221_barrel_shifter_line72 = {tmp220_barrel_shifter_line72};
    assign tmp222_barrel_shifter_line72 = tmp219_barrel_shifter_line72 | tmp221_barrel_shifter_line72;
    assign tmp223_barrel_shifter_line72 = {tmp216_barrel_shifter_line72[3], tmp216_barrel_shifter_line72[2]};
    assign tmp224_barrel_shifter_line72 = {tmp223_barrel_shifter_line72[0]};
    assign tmp225_barrel_shifter_line72 = {tmp224_barrel_shifter_line72};
    assign tmp226_barrel_shifter_line72 = {tmp223_barrel_shifter_line72[1]};
    assign tmp227_barrel_shifter_line72 = {tmp226_barrel_shifter_line72};
    assign tmp228_barrel_shifter_line72 = tmp225_barrel_shifter_line72 | tmp227_barrel_shifter_line72;
    assign tmp229_barrel_shifter_line72 = tmp222_barrel_shifter_line72 | tmp228_barrel_shifter_line72;
    assign tmp230_barrel_shifter_line72 = tmp215_barrel_shifter_line72 | tmp229_barrel_shifter_line72;
    assign tmp231_barrel_shifter_line72 = {tmp200_barrel_shifter_line72[15], tmp200_barrel_shifter_line72[14], tmp200_barrel_shifter_line72[13], tmp200_barrel_shifter_line72[12], tmp200_barrel_shifter_line72[11], tmp200_barrel_shifter_line72[10], tmp200_barrel_shifter_line72[9], tmp200_barrel_shifter_line72[8]};
    assign tmp232_barrel_shifter_line72 = {tmp231_barrel_shifter_line72[3], tmp231_barrel_shifter_line72[2], tmp231_barrel_shifter_line72[1], tmp231_barrel_shifter_line72[0]};
    assign tmp233_barrel_shifter_line72 = {tmp232_barrel_shifter_line72[1], tmp232_barrel_shifter_line72[0]};
    assign tmp234_barrel_shifter_line72 = {tmp233_barrel_shifter_line72[0]};
    assign tmp235_barrel_shifter_line72 = {tmp234_barrel_shifter_line72};
    assign tmp236_barrel_shifter_line72 = {tmp233_barrel_shifter_line72[1]};
    assign tmp237_barrel_shifter_line72 = {tmp236_barrel_shifter_line72};
    assign tmp238_barrel_shifter_line72 = tmp235_barrel_shifter_line72 | tmp237_barrel_shifter_line72;
    assign tmp239_barrel_shifter_line72 = {tmp232_barrel_shifter_line72[3], tmp232_barrel_shifter_line72[2]};
    assign tmp240_barrel_shifter_line72 = {tmp239_barrel_shifter_line72[0]};
    assign tmp241_barrel_shifter_line72 = {tmp240_barrel_shifter_line72};
    assign tmp242_barrel_shifter_line72 = {tmp239_barrel_shifter_line72[1]};
    assign tmp243_barrel_shifter_line72 = {tmp242_barrel_shifter_line72};
    assign tmp244_barrel_shifter_line72 = tmp241_barrel_shifter_line72 | tmp243_barrel_shifter_line72;
    assign tmp245_barrel_shifter_line72 = tmp238_barrel_shifter_line72 | tmp244_barrel_shifter_line72;
    assign tmp246_barrel_shifter_line72 = {tmp231_barrel_shifter_line72[7], tmp231_barrel_shifter_line72[6], tmp231_barrel_shifter_line72[5], tmp231_barrel_shifter_line72[4]};
    assign tmp247_barrel_shifter_line72 = {tmp246_barrel_shifter_line72[1], tmp246_barrel_shifter_line72[0]};
    assign tmp248_barrel_shifter_line72 = {tmp247_barrel_shifter_line72[0]};
    assign tmp249_barrel_shifter_line72 = {tmp248_barrel_shifter_line72};
    assign tmp250_barrel_shifter_line72 = {tmp247_barrel_shifter_line72[1]};
    assign tmp251_barrel_shifter_line72 = {tmp250_barrel_shifter_line72};
    assign tmp252_barrel_shifter_line72 = tmp249_barrel_shifter_line72 | tmp251_barrel_shifter_line72;
    assign tmp253_barrel_shifter_line72 = {tmp246_barrel_shifter_line72[3], tmp246_barrel_shifter_line72[2]};
    assign tmp254_barrel_shifter_line72 = {tmp253_barrel_shifter_line72[0]};
    assign tmp255_barrel_shifter_line72 = {tmp254_barrel_shifter_line72};
    assign tmp256_barrel_shifter_line72 = {tmp253_barrel_shifter_line72[1]};
    assign tmp257_barrel_shifter_line72 = {tmp256_barrel_shifter_line72};
    assign tmp258_barrel_shifter_line72 = tmp255_barrel_shifter_line72 | tmp257_barrel_shifter_line72;
    assign tmp259_barrel_shifter_line72 = tmp252_barrel_shifter_line72 | tmp258_barrel_shifter_line72;
    assign tmp260_barrel_shifter_line72 = tmp245_barrel_shifter_line72 | tmp259_barrel_shifter_line72;
    assign tmp261_barrel_shifter_line72 = tmp230_barrel_shifter_line72 | tmp260_barrel_shifter_line72;
    assign tmp262_barrel_shifter_line72 = {shift_off_32[31], shift_off_32[30], shift_off_32[29], shift_off_32[28], shift_off_32[27], shift_off_32[26], shift_off_32[25], shift_off_32[24], shift_off_32[23], shift_off_32[22], shift_off_32[21], shift_off_32[20], shift_off_32[19], shift_off_32[18], shift_off_32[17], shift_off_32[16]};
    assign tmp263_barrel_shifter_line72 = {tmp262_barrel_shifter_line72[7], tmp262_barrel_shifter_line72[6], tmp262_barrel_shifter_line72[5], tmp262_barrel_shifter_line72[4], tmp262_barrel_shifter_line72[3], tmp262_barrel_shifter_line72[2], tmp262_barrel_shifter_line72[1], tmp262_barrel_shifter_line72[0]};
    assign tmp264_barrel_shifter_line72 = {tmp263_barrel_shifter_line72[3], tmp263_barrel_shifter_line72[2], tmp263_barrel_shifter_line72[1], tmp263_barrel_shifter_line72[0]};
    assign tmp265_barrel_shifter_line72 = {tmp264_barrel_shifter_line72[1], tmp264_barrel_shifter_line72[0]};
    assign tmp266_barrel_shifter_line72 = {tmp265_barrel_shifter_line72[0]};
    assign tmp267_barrel_shifter_line72 = {tmp266_barrel_shifter_line72};
    assign tmp268_barrel_shifter_line72 = {tmp265_barrel_shifter_line72[1]};
    assign tmp269_barrel_shifter_line72 = {tmp268_barrel_shifter_line72};
    assign tmp270_barrel_shifter_line72 = tmp267_barrel_shifter_line72 | tmp269_barrel_shifter_line72;
    assign tmp271_barrel_shifter_line72 = {tmp264_barrel_shifter_line72[3], tmp264_barrel_shifter_line72[2]};
    assign tmp272_barrel_shifter_line72 = {tmp271_barrel_shifter_line72[0]};
    assign tmp273_barrel_shifter_line72 = {tmp272_barrel_shifter_line72};
    assign tmp274_barrel_shifter_line72 = {tmp271_barrel_shifter_line72[1]};
    assign tmp275_barrel_shifter_line72 = {tmp274_barrel_shifter_line72};
    assign tmp276_barrel_shifter_line72 = tmp273_barrel_shifter_line72 | tmp275_barrel_shifter_line72;
    assign tmp277_barrel_shifter_line72 = tmp270_barrel_shifter_line72 | tmp276_barrel_shifter_line72;
    assign tmp278_barrel_shifter_line72 = {tmp263_barrel_shifter_line72[7], tmp263_barrel_shifter_line72[6], tmp263_barrel_shifter_line72[5], tmp263_barrel_shifter_line72[4]};
    assign tmp279_barrel_shifter_line72 = {tmp278_barrel_shifter_line72[1], tmp278_barrel_shifter_line72[0]};
    assign tmp280_barrel_shifter_line72 = {tmp279_barrel_shifter_line72[0]};
    assign tmp281_barrel_shifter_line72 = {tmp280_barrel_shifter_line72};
    assign tmp282_barrel_shifter_line72 = {tmp279_barrel_shifter_line72[1]};
    assign tmp283_barrel_shifter_line72 = {tmp282_barrel_shifter_line72};
    assign tmp284_barrel_shifter_line72 = tmp281_barrel_shifter_line72 | tmp283_barrel_shifter_line72;
    assign tmp285_barrel_shifter_line72 = {tmp278_barrel_shifter_line72[3], tmp278_barrel_shifter_line72[2]};
    assign tmp286_barrel_shifter_line72 = {tmp285_barrel_shifter_line72[0]};
    assign tmp287_barrel_shifter_line72 = {tmp286_barrel_shifter_line72};
    assign tmp288_barrel_shifter_line72 = {tmp285_barrel_shifter_line72[1]};
    assign tmp289_barrel_shifter_line72 = {tmp288_barrel_shifter_line72};
    assign tmp290_barrel_shifter_line72 = tmp287_barrel_shifter_line72 | tmp289_barrel_shifter_line72;
    assign tmp291_barrel_shifter_line72 = tmp284_barrel_shifter_line72 | tmp290_barrel_shifter_line72;
    assign tmp292_barrel_shifter_line72 = tmp277_barrel_shifter_line72 | tmp291_barrel_shifter_line72;
    assign tmp293_barrel_shifter_line72 = {tmp262_barrel_shifter_line72[15], tmp262_barrel_shifter_line72[14], tmp262_barrel_shifter_line72[13], tmp262_barrel_shifter_line72[12], tmp262_barrel_shifter_line72[11], tmp262_barrel_shifter_line72[10], tmp262_barrel_shifter_line72[9], tmp262_barrel_shifter_line72[8]};
    assign tmp294_barrel_shifter_line72 = {tmp293_barrel_shifter_line72[3], tmp293_barrel_shifter_line72[2], tmp293_barrel_shifter_line72[1], tmp293_barrel_shifter_line72[0]};
    assign tmp295_barrel_shifter_line72 = {tmp294_barrel_shifter_line72[1], tmp294_barrel_shifter_line72[0]};
    assign tmp296_barrel_shifter_line72 = {tmp295_barrel_shifter_line72[0]};
    assign tmp297_barrel_shifter_line72 = {tmp296_barrel_shifter_line72};
    assign tmp298_barrel_shifter_line72 = {tmp295_barrel_shifter_line72[1]};
    assign tmp299_barrel_shifter_line72 = {tmp298_barrel_shifter_line72};
    assign tmp300_barrel_shifter_line72 = tmp297_barrel_shifter_line72 | tmp299_barrel_shifter_line72;
    assign tmp301_barrel_shifter_line72 = {tmp294_barrel_shifter_line72[3], tmp294_barrel_shifter_line72[2]};
    assign tmp302_barrel_shifter_line72 = {tmp301_barrel_shifter_line72[0]};
    assign tmp303_barrel_shifter_line72 = {tmp302_barrel_shifter_line72};
    assign tmp304_barrel_shifter_line72 = {tmp301_barrel_shifter_line72[1]};
    assign tmp305_barrel_shifter_line72 = {tmp304_barrel_shifter_line72};
    assign tmp306_barrel_shifter_line72 = tmp303_barrel_shifter_line72 | tmp305_barrel_shifter_line72;
    assign tmp307_barrel_shifter_line72 = tmp300_barrel_shifter_line72 | tmp306_barrel_shifter_line72;
    assign tmp308_barrel_shifter_line72 = {tmp293_barrel_shifter_line72[7], tmp293_barrel_shifter_line72[6], tmp293_barrel_shifter_line72[5], tmp293_barrel_shifter_line72[4]};
    assign tmp309_barrel_shifter_line72 = {tmp308_barrel_shifter_line72[1], tmp308_barrel_shifter_line72[0]};
    assign tmp310_barrel_shifter_line72 = {tmp309_barrel_shifter_line72[0]};
    assign tmp311_barrel_shifter_line72 = {tmp310_barrel_shifter_line72};
    assign tmp312_barrel_shifter_line72 = {tmp309_barrel_shifter_line72[1]};
    assign tmp313_barrel_shifter_line72 = {tmp312_barrel_shifter_line72};
    assign tmp314_barrel_shifter_line72 = tmp311_barrel_shifter_line72 | tmp313_barrel_shifter_line72;
    assign tmp315_barrel_shifter_line72 = {tmp308_barrel_shifter_line72[3], tmp308_barrel_shifter_line72[2]};
    assign tmp316_barrel_shifter_line72 = {tmp315_barrel_shifter_line72[0]};
    assign tmp317_barrel_shifter_line72 = {tmp316_barrel_shifter_line72};
    assign tmp318_barrel_shifter_line72 = {tmp315_barrel_shifter_line72[1]};
    assign tmp319_barrel_shifter_line72 = {tmp318_barrel_shifter_line72};
    assign tmp320_barrel_shifter_line72 = tmp317_barrel_shifter_line72 | tmp319_barrel_shifter_line72;
    assign tmp321_barrel_shifter_line72 = tmp314_barrel_shifter_line72 | tmp320_barrel_shifter_line72;
    assign tmp322_barrel_shifter_line72 = tmp307_barrel_shifter_line72 | tmp321_barrel_shifter_line72;
    assign tmp323_barrel_shifter_line72 = tmp292_barrel_shifter_line72 | tmp322_barrel_shifter_line72;
    assign tmp324_barrel_shifter_line72 = tmp261_barrel_shifter_line72 | tmp323_barrel_shifter_line72;
    assign tmp325_barrel_shifter_line72 = {shift_off_16[7], shift_off_16[6], shift_off_16[5], shift_off_16[4], shift_off_16[3], shift_off_16[2], shift_off_16[1], shift_off_16[0]};
    assign tmp326_barrel_shifter_line72 = {tmp325_barrel_shifter_line72[3], tmp325_barrel_shifter_line72[2], tmp325_barrel_shifter_line72[1], tmp325_barrel_shifter_line72[0]};
    assign tmp327_barrel_shifter_line72 = {tmp326_barrel_shifter_line72[1], tmp326_barrel_shifter_line72[0]};
    assign tmp328_barrel_shifter_line72 = {tmp327_barrel_shifter_line72[0]};
    assign tmp329_barrel_shifter_line72 = {tmp328_barrel_shifter_line72};
    assign tmp330_barrel_shifter_line72 = {tmp327_barrel_shifter_line72[1]};
    assign tmp331_barrel_shifter_line72 = {tmp330_barrel_shifter_line72};
    assign tmp332_barrel_shifter_line72 = tmp329_barrel_shifter_line72 | tmp331_barrel_shifter_line72;
    assign tmp333_barrel_shifter_line72 = {tmp326_barrel_shifter_line72[3], tmp326_barrel_shifter_line72[2]};
    assign tmp334_barrel_shifter_line72 = {tmp333_barrel_shifter_line72[0]};
    assign tmp335_barrel_shifter_line72 = {tmp334_barrel_shifter_line72};
    assign tmp336_barrel_shifter_line72 = {tmp333_barrel_shifter_line72[1]};
    assign tmp337_barrel_shifter_line72 = {tmp336_barrel_shifter_line72};
    assign tmp338_barrel_shifter_line72 = tmp335_barrel_shifter_line72 | tmp337_barrel_shifter_line72;
    assign tmp339_barrel_shifter_line72 = tmp332_barrel_shifter_line72 | tmp338_barrel_shifter_line72;
    assign tmp340_barrel_shifter_line72 = {tmp325_barrel_shifter_line72[7], tmp325_barrel_shifter_line72[6], tmp325_barrel_shifter_line72[5], tmp325_barrel_shifter_line72[4]};
    assign tmp341_barrel_shifter_line72 = {tmp340_barrel_shifter_line72[1], tmp340_barrel_shifter_line72[0]};
    assign tmp342_barrel_shifter_line72 = {tmp341_barrel_shifter_line72[0]};
    assign tmp343_barrel_shifter_line72 = {tmp342_barrel_shifter_line72};
    assign tmp344_barrel_shifter_line72 = {tmp341_barrel_shifter_line72[1]};
    assign tmp345_barrel_shifter_line72 = {tmp344_barrel_shifter_line72};
    assign tmp346_barrel_shifter_line72 = tmp343_barrel_shifter_line72 | tmp345_barrel_shifter_line72;
    assign tmp347_barrel_shifter_line72 = {tmp340_barrel_shifter_line72[3], tmp340_barrel_shifter_line72[2]};
    assign tmp348_barrel_shifter_line72 = {tmp347_barrel_shifter_line72[0]};
    assign tmp349_barrel_shifter_line72 = {tmp348_barrel_shifter_line72};
    assign tmp350_barrel_shifter_line72 = {tmp347_barrel_shifter_line72[1]};
    assign tmp351_barrel_shifter_line72 = {tmp350_barrel_shifter_line72};
    assign tmp352_barrel_shifter_line72 = tmp349_barrel_shifter_line72 | tmp351_barrel_shifter_line72;
    assign tmp353_barrel_shifter_line72 = tmp346_barrel_shifter_line72 | tmp352_barrel_shifter_line72;
    assign tmp354_barrel_shifter_line72 = tmp339_barrel_shifter_line72 | tmp353_barrel_shifter_line72;
    assign tmp355_barrel_shifter_line72 = {shift_off_16[15], shift_off_16[14], shift_off_16[13], shift_off_16[12], shift_off_16[11], shift_off_16[10], shift_off_16[9], shift_off_16[8]};
    assign tmp356_barrel_shifter_line72 = {tmp355_barrel_shifter_line72[3], tmp355_barrel_shifter_line72[2], tmp355_barrel_shifter_line72[1], tmp355_barrel_shifter_line72[0]};
    assign tmp357_barrel_shifter_line72 = {tmp356_barrel_shifter_line72[1], tmp356_barrel_shifter_line72[0]};
    assign tmp358_barrel_shifter_line72 = {tmp357_barrel_shifter_line72[0]};
    assign tmp359_barrel_shifter_line72 = {tmp358_barrel_shifter_line72};
    assign tmp360_barrel_shifter_line72 = {tmp357_barrel_shifter_line72[1]};
    assign tmp361_barrel_shifter_line72 = {tmp360_barrel_shifter_line72};
    assign tmp362_barrel_shifter_line72 = tmp359_barrel_shifter_line72 | tmp361_barrel_shifter_line72;
    assign tmp363_barrel_shifter_line72 = {tmp356_barrel_shifter_line72[3], tmp356_barrel_shifter_line72[2]};
    assign tmp364_barrel_shifter_line72 = {tmp363_barrel_shifter_line72[0]};
    assign tmp365_barrel_shifter_line72 = {tmp364_barrel_shifter_line72};
    assign tmp366_barrel_shifter_line72 = {tmp363_barrel_shifter_line72[1]};
    assign tmp367_barrel_shifter_line72 = {tmp366_barrel_shifter_line72};
    assign tmp368_barrel_shifter_line72 = tmp365_barrel_shifter_line72 | tmp367_barrel_shifter_line72;
    assign tmp369_barrel_shifter_line72 = tmp362_barrel_shifter_line72 | tmp368_barrel_shifter_line72;
    assign tmp370_barrel_shifter_line72 = {tmp355_barrel_shifter_line72[7], tmp355_barrel_shifter_line72[6], tmp355_barrel_shifter_line72[5], tmp355_barrel_shifter_line72[4]};
    assign tmp371_barrel_shifter_line72 = {tmp370_barrel_shifter_line72[1], tmp370_barrel_shifter_line72[0]};
    assign tmp372_barrel_shifter_line72 = {tmp371_barrel_shifter_line72[0]};
    assign tmp373_barrel_shifter_line72 = {tmp372_barrel_shifter_line72};
    assign tmp374_barrel_shifter_line72 = {tmp371_barrel_shifter_line72[1]};
    assign tmp375_barrel_shifter_line72 = {tmp374_barrel_shifter_line72};
    assign tmp376_barrel_shifter_line72 = tmp373_barrel_shifter_line72 | tmp375_barrel_shifter_line72;
    assign tmp377_barrel_shifter_line72 = {tmp370_barrel_shifter_line72[3], tmp370_barrel_shifter_line72[2]};
    assign tmp378_barrel_shifter_line72 = {tmp377_barrel_shifter_line72[0]};
    assign tmp379_barrel_shifter_line72 = {tmp378_barrel_shifter_line72};
    assign tmp380_barrel_shifter_line72 = {tmp377_barrel_shifter_line72[1]};
    assign tmp381_barrel_shifter_line72 = {tmp380_barrel_shifter_line72};
    assign tmp382_barrel_shifter_line72 = tmp379_barrel_shifter_line72 | tmp381_barrel_shifter_line72;
    assign tmp383_barrel_shifter_line72 = tmp376_barrel_shifter_line72 | tmp382_barrel_shifter_line72;
    assign tmp384_barrel_shifter_line72 = tmp369_barrel_shifter_line72 | tmp383_barrel_shifter_line72;
    assign tmp385_barrel_shifter_line72 = tmp354_barrel_shifter_line72 | tmp384_barrel_shifter_line72;
    assign tmp386_barrel_shifter_line72 = tmp324_barrel_shifter_line72 | tmp385_barrel_shifter_line72;
    assign tmp387_barrel_shifter_line72 = {shift_off_8[3], shift_off_8[2], shift_off_8[1], shift_off_8[0]};
    assign tmp388_barrel_shifter_line72 = {tmp387_barrel_shifter_line72[1], tmp387_barrel_shifter_line72[0]};
    assign tmp389_barrel_shifter_line72 = {tmp388_barrel_shifter_line72[0]};
    assign tmp390_barrel_shifter_line72 = {tmp389_barrel_shifter_line72};
    assign tmp391_barrel_shifter_line72 = {tmp388_barrel_shifter_line72[1]};
    assign tmp392_barrel_shifter_line72 = {tmp391_barrel_shifter_line72};
    assign tmp393_barrel_shifter_line72 = tmp390_barrel_shifter_line72 | tmp392_barrel_shifter_line72;
    assign tmp394_barrel_shifter_line72 = {tmp387_barrel_shifter_line72[3], tmp387_barrel_shifter_line72[2]};
    assign tmp395_barrel_shifter_line72 = {tmp394_barrel_shifter_line72[0]};
    assign tmp396_barrel_shifter_line72 = {tmp395_barrel_shifter_line72};
    assign tmp397_barrel_shifter_line72 = {tmp394_barrel_shifter_line72[1]};
    assign tmp398_barrel_shifter_line72 = {tmp397_barrel_shifter_line72};
    assign tmp399_barrel_shifter_line72 = tmp396_barrel_shifter_line72 | tmp398_barrel_shifter_line72;
    assign tmp400_barrel_shifter_line72 = tmp393_barrel_shifter_line72 | tmp399_barrel_shifter_line72;
    assign tmp401_barrel_shifter_line72 = {shift_off_8[7], shift_off_8[6], shift_off_8[5], shift_off_8[4]};
    assign tmp402_barrel_shifter_line72 = {tmp401_barrel_shifter_line72[1], tmp401_barrel_shifter_line72[0]};
    assign tmp403_barrel_shifter_line72 = {tmp402_barrel_shifter_line72[0]};
    assign tmp404_barrel_shifter_line72 = {tmp403_barrel_shifter_line72};
    assign tmp405_barrel_shifter_line72 = {tmp402_barrel_shifter_line72[1]};
    assign tmp406_barrel_shifter_line72 = {tmp405_barrel_shifter_line72};
    assign tmp407_barrel_shifter_line72 = tmp404_barrel_shifter_line72 | tmp406_barrel_shifter_line72;
    assign tmp408_barrel_shifter_line72 = {tmp401_barrel_shifter_line72[3], tmp401_barrel_shifter_line72[2]};
    assign tmp409_barrel_shifter_line72 = {tmp408_barrel_shifter_line72[0]};
    assign tmp410_barrel_shifter_line72 = {tmp409_barrel_shifter_line72};
    assign tmp411_barrel_shifter_line72 = {tmp408_barrel_shifter_line72[1]};
    assign tmp412_barrel_shifter_line72 = {tmp411_barrel_shifter_line72};
    assign tmp413_barrel_shifter_line72 = tmp410_barrel_shifter_line72 | tmp412_barrel_shifter_line72;
    assign tmp414_barrel_shifter_line72 = tmp407_barrel_shifter_line72 | tmp413_barrel_shifter_line72;
    assign tmp415_barrel_shifter_line72 = tmp400_barrel_shifter_line72 | tmp414_barrel_shifter_line72;
    assign tmp416_barrel_shifter_line72 = tmp386_barrel_shifter_line72 | tmp415_barrel_shifter_line72;
    assign tmp417_barrel_shifter_line72 = {shift_off_4[1], shift_off_4[0]};
    assign tmp418_barrel_shifter_line72 = {tmp417_barrel_shifter_line72[0]};
    assign tmp419_barrel_shifter_line72 = {tmp418_barrel_shifter_line72};
    assign tmp420_barrel_shifter_line72 = {tmp417_barrel_shifter_line72[1]};
    assign tmp421_barrel_shifter_line72 = {tmp420_barrel_shifter_line72};
    assign tmp422_barrel_shifter_line72 = tmp419_barrel_shifter_line72 | tmp421_barrel_shifter_line72;
    assign tmp423_barrel_shifter_line72 = {shift_off_4[3], shift_off_4[2]};
    assign tmp424_barrel_shifter_line72 = {tmp423_barrel_shifter_line72[0]};
    assign tmp425_barrel_shifter_line72 = {tmp424_barrel_shifter_line72};
    assign tmp426_barrel_shifter_line72 = {tmp423_barrel_shifter_line72[1]};
    assign tmp427_barrel_shifter_line72 = {tmp426_barrel_shifter_line72};
    assign tmp428_barrel_shifter_line72 = tmp425_barrel_shifter_line72 | tmp427_barrel_shifter_line72;
    assign tmp429_barrel_shifter_line72 = tmp422_barrel_shifter_line72 | tmp428_barrel_shifter_line72;
    assign tmp430_barrel_shifter_line72 = tmp416_barrel_shifter_line72 | tmp429_barrel_shifter_line72;
    assign tmp431_barrel_shifter_line72 = {shift_off_2[0]};
    assign tmp432_barrel_shifter_line72 = {tmp431_barrel_shifter_line72};
    assign tmp433_barrel_shifter_line72 = {shift_off_2[1]};
    assign tmp434_barrel_shifter_line72 = {tmp433_barrel_shifter_line72};
    assign tmp435_barrel_shifter_line72 = tmp432_barrel_shifter_line72 | tmp434_barrel_shifter_line72;
    assign tmp436_barrel_shifter_line72 = tmp430_barrel_shifter_line72 | tmp435_barrel_shifter_line72;
    assign tmp437_barrel_shifter_line72 = {shift_off_1};
    assign tmp438_barrel_shifter_line72 = tmp436_barrel_shifter_line72 | tmp437_barrel_shifter_line72;

endmodule
